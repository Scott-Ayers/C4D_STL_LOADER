MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ��P�یP�یP�ی�2�Q�ی]��N�ی]�:��ی]�;���ی�m�S�یP�ڌ�ی�:�J�ی��Q�ی��Q�یRichP�ی                PE  L P�Z        � !  "  f     �.                               �         @                   p� [  � (                              �  �_ 8                           8 @             �                          .textbss�                        �  �.text   y!     "                   `.rdata  �\  P  ^  &             @  @.data   �_   �  2   �             @  �.idata  �        �             @  @.reloc  ��      �   �             @  B                                                                                                                                                                                                                                                                                                        ������ �a� ��� 駟 �2� �- �� �� ��Z �9B �4� �Oj �5 ��X �> �~ ��� ��p �� �� �M �]� �s �S�
 �.� 鹓 �, �?� �
� �e ��� �o	 �F 鑥 �� ��o �� �� �Lj �c� �N9 �Yt ��� �_a
 銌 �K ��@ �  �V� ��' �L@ �ǖ �
 �]� � �% ��~ ��� �D�  ��� 骳 �uW ��b	 � �M �! �v	 �G �"� �=� �X� �se
 �~� �9� 餢 �� ��� �� ��� �[� ��I	 �1� �l �� �" ��	 �� �## �6 �ə �� �oz �: ��) ��� �;n �v�	 �q� ��� �w� �> 靼 � 飤 �� �i �� �� ��  �EN ��� �s �6j �a� ��$ �7 �n �� ��� �3n �� �� �� �!
 �. �5� 鰀 �[� �v� 鑶 �( �1 ��� �m� �H� �� ��� ��� �h �_�  �J� �U �L �{ 鶆 �� �� �� �R9 �]� ��R ��� ��u
 �)�	 �t� ��f �
�	 �u� �`b �k �FG �o �� �7 �* �c �& �c� �� � �D� ��	 �e �G �� �t �� �1 �Hg �7G �� �}� �f �c� ��
 �i% �d �� ��c	 ��F ��� ���  ��{ �A� �f �g�
 �Bs ��� ��� �#0 �� ��C �& �  �2
 �R � � ��g �ƈ ��  �\S
 �$
 �
g �}� �H �n �r �	� �� �/� �� �� �  髱 ��  �g
 鼅 ��	 �, �� ��� �? ��� �6 �$Q �� �) ��� �`G ��� �F ��0 �* ��
 ��� �T �� ���
 �9 �y �f �� �
" �� �0� ��� �� �aU �M � �b� ��l �(S ��� �pe �	u �V ��T � �e� �p� �� �v�  �� 鼬 ��� �R� ��P �X ��d � �i& � �?"
 �z� �5� �P� �ˎ	 �[ �' ��  �W' �"� �� ��P �c	 �� �Is �d �d ��E �r �@C �� �� 遤 ���  �g� �� �� �; ��6 �^s �I�  �d� �?� ��/
 �%� �p� � �F] �q: ��	 �w� ��� �-� �8s �3 �� �y� �� ��� �j�	 ��� ��S �[" �G
 ��	 ��b �w� ��� �= ��s �3a �.� �)P �� �?d �D
 ��p �`� 雟 �V]	 �� �l �g� 钑 �}� �� ��7 �.V ��L 鄤 �/d �� � �p� � ��� �X �LW ��� �_	 �Ͷ �� �sf �e �9� �� �  �� 酸 ��y �j �� �Q� �g ��' �r�	 �� �hj ���  ��
 ��* �d( �� �g �e
 � & � �6� �� �L� �'a ��_ �R �hn
 �cF �>6 �� ��� 韨 �J8 鵩 �p� ��n ��� 鑧 �<� ��' ��/ ��	 �b �C� �� �� ��� ��� ��� ��j ��� � ��� �[ �L� �# �G �m �(�  �3S ��=	 �)�  ��E �2 ��b ���  �P; ��� �V� �Q� ��� �w �B7	 ��V
 �O ��F � ��B �4x � �*| �U�  �PN ��c �l �j �,i �w� �x �c �Nb �Ӌ	 ��� �i� 鴯 ��� �� ��4 �P& �O �fg �qe � �w4 ���
 �}� �0 �3� �^� �I6	 ��l ���  �3 �5 �@+ �[4 ��� �_ �, ��v ��x ��	 ��? �s� �^� ��H �a �?
 �J� �ui
 �� ��� ��  �� �; �W� �bO
 �� �] �o ��� �y� �$� 韌 ��q �� �  �C �f[	 �� �<� �U ��A �}� �H� �t �~� �� �e �� �� 饐 �@� �� ��_ ��� �\� �e ��� �-� �  ��[	 �! �	 ��4 ���
 ��� �5~ �@� ��`
 �� �F �L` ��� ��� �h �x ���  ��	 �	�  鴩 鿵  麩 �u� ��C �$ �fC �� �� �gC �R� ��K
 ��  �3 �.�	 �y� ��� 鏰 � ��� � ��% � ��< ��� ��� �R�
 �I
 �< �� � �i	 �İ � �ʊ �� �� ��& �6� �a�
 ��� ��7 �R3 � �H� �- �� �y� �46 �O� �*� �el ��I �{� �A �a� �� �G
 �� ��� 阯 �S^ � �	�  ��� �� �:T �� �  ��Q �F �A �L� � �RZ	 �$
 �7 �� �^w �yJ ��� �_� �� �� � �6 � �Q� �|! ��_ �BL 靉 �_ �= �N � �4, �� ��] 鵳 �P� �, �&k ��J �� � �bI ��r �( �#� � �	� �Tv �/ �� �� �p> �K�	 �V �QV ���  ��� ��� � 阊 �CN ��
 �)� �$� �O �: �� �p� �� ��� 遠	 �< ��� ��  �m� �� 铕 ��d �)� ��: ��O ��� ��3 ��J ��� �F� ��� �6 �W� �B �M> �� �C� �.M	 �� �� ���  �Jc �] �p= �+- �f�  ��� �l� ��� ���
 �-n �( �} �.� �)� �; ��" �� �
 �� �� �� ��b �< �g �B�
 �M ��  �8� 龫 �	� ��	 ��@	 ��\ �%l �j �{�
 ��  �q� �� �G 鲟 ��	 �/ � �� �i� �D� �_�	 �! ��� �" �Kt �o �X	 �<� �� �B�
 ��	 �(� � �N� �� �t� �' ��[ �uo �`�  �[G
 �V �a  �| �'� �� �< �8� �3I �F �9� ��[ � �0 �� �Z � �6� 顫 ���  �7� ��^ �mf
 �x� �C �� ��? �$ �o� ��  �U� �P �K� �H
 �1� �� ��Y �i �-l �H[ ���
 �C
 �I� �� ��	 �ک 镗 �� �+� �f �� ��� �'� �Q �-�	 �[ �a
 龡 � �DW �/? �� �e� 須 �V	 鶠 �QE � ��
 ��L �m ��v �� �N: �� �4 鏰 �z> �U/ � T	 �۩ ��W �� ��� � �tZ �z �(� �� �6 �i �D�	 �� �*� �1u �� �+  ��* �!H �\�  �'� 鲦
 �y �Ȋ �F	 �� �"�	 �ı  �OO
 �z� �u � T	 �;� �� �� �: ��� �� ���	 �� �� 鎡 �� �� �0
 �:� �U� �g� �;o	 �� �1�  �L� �`
 �2�  �} � 郰 �N� ��1 ��" �& ��	 鵪 �P �k �V� ��2 鬀 ��@ �"� �� �(� 铖 �~� �I� �$� �� �� � � 雯 �a ��o ��
 ���	 �2� ��F ��� �� �n6 �i� �: �O� 麮 �E	 �`� �� �A �� 鬕 釔 �B� �	 �X� �c� �n�  �٤
 ���  ��c �� �� �P� �( �v� �� � �G] �B  �=_
 �� �C� �e ��k	 �� 鿨 �: �E�  ��O �� ��{ �q� ��! �� �
 �� �Xv ��. �� ��) �� ��	 ��� 酄 �0*	 �k�	 ��� �Q� ��c 鷀	 �B: �m 阾
 �c�	 �N	 �	� �D �� ��h �յ	 �`
 � �� �& � 鷘 针 �m� �h� �s0 �^�
 �� ��  �O/ �JS ��� 頝 ��& ��� �1� ��� �Ǫ � �� �� �� ��� ��� �D� �� 銨 ��
 頬 髞 �� ��5 �\	 �� �B� �� ��� �� ��� ��f �4  �O� 麋 �u� ��� 雷 � �� �<8 �w� �! ��� �� �s� ��- �	� �� � ��; ��  ��	 ��� ��� �K �L� �� �"�  ��
 �� �� � �9�	 �t ��> �� �Ey �? ��| ��s ��
 �,n �u 邋 �]7 �، �cO �~� ��� �M �o �j� �� � � ��� �&N �A �Z �י 额 �=o ��8 �s �N! �0 �ԋ �� �J2 � �p �[L 醔 �!1 �L�
 �w �" �]�  �?
 �c �F �9& ��  �/�  �� �e
 ��� ��	 ��n �a| �L8 �W( �r� �n ��� �s� �> �	� �T� �?� �ʵ ��k	 �Ps �� �F� � � �Wn �R �=U
 ��� �SY �^y �i �  ��  �J� �I � � �kL	 ���  �Ae ��  �� ��� ���  �� �3 �N� � ��� ��	 �j� �s �� �o �� �1W �D �p �rX
 �S	 ��m ��� �P �y �4B �O� �j�
 �E� ��� � �� �a\ �L�	 �g	 �r  �� �. �s� �. ��  ��
 �i� ��' �E�
 �p
 �{� �v� �) � �� �ҥ �-�  ��� �3B �n �9 �d� �} ��1 �k �B �� �  鑵 �� �w� � ��� �8F � �K	 �� �d� �Χ �ʙ �E �P� ��V
 �։
 �� �� �'�  �2� �� �8 ��
 �NG ��� �� �� 隹 �� �% �{� ��p ��/ �|= �� �B� �aR �
 �z �' �	X
 � �� �Z�
 �OQ �� �; ��Q
 遂 �p �
 �R
 靋 �I	 ��, �� �� �T  �B �*� �� � �{z ��� �QC �� �7�  �r� ���
 �� �| �Q ��� �� ��� ���  �D 鐱 ��: �	 �ad ���  �cQ �R#	 �Y ���  ��
 �^ �y �� �/� �z� �5U �p� �� � �a� ��	 �} �"�  � �H4 ��A ��� ��� ��t �� �� �J	 � 1 ��t ��� �!� 鼭	 � �2O � � �� �.�  �ً �l �O7 ��� �E�  ��	 ��� �Ư ��� � �R �2 �- �8� ��T �� �ij �: �o� �Z �� � [ �[�	 �,	 �! ��e �~ �R� � ��4 �3t �^� �I4 �� �� ��N � 逨 �{� 鶗	 ��� �� �w� � �]� �(� ���  �V� �	� �Ę � �J� ��� � � �� ���  ��? �q �= �"� �� �(U
 ��� � �)2 �N 韰 �� �X ���  �� �� �� �lz � ��-	 �� �h1 ���	 �^� �y.	 �� � �� ��M �p{ �� �C �� �,� �w �� ��> �H	 � �! �)�
 ��{ �_� �z+ �) 鰓 雄 �jM ��m �<�  �7 �W
 �-� �� �� �� �Q �� ��  �I ��' �0 �{� ��� �1� �&
 �7� � ��| ��� �C� 龍 �y� �ԅ �L �ʞ
 �L � | ��� �&8
 ��� �<�
 �'7 � � �� �CK ��  ��j �T� 韁 � �_L �� �ہ �v� �o ���  �� ��  �M�	 �� ��l ��R ��
 �4] � �ZR �E� �л
 �;�	 � �a� �8 �v �� ��\ �H� �#} �� 陯 餫 �� �� ���
 ���
 �8
 �V�
 鑫 �� �W� �� �� �� ��� �j �I� �t  �_ �:^ ���  ���  �[�  �&� �� �ܜ �� ��� �� �� ��
 ��� �IG �tv ��*	 �� �%~ �� �[ �ր ��w �n �B �җ ��
 �� �� �� ���
 �D �?x �:Q �� �� �� �L 顜	 �<� �� ��� �iL �$ �S  �΀	 �	� � 鯫 �j� �%�
 �p �{�	 �&& �1F	 �/ �UJ ��� �?
 ��	 飩 ��  �� �dI �o�  �
 ��  �� ��" �/ �!R �| �w� �� �m� �X�  ��� �>r ��
 �) �/� ��3
 �� �  �8
 �6�  � � �g7 �b� �� �X� �÷  �� 驹  鴔 ��� �u �59 � � �+� � ��M
 �L� �g# ��I �� �� ��< �� �t � ��
 �: ��P �� �� �v�
 �AE
 �<� �z �? �O �� �3Q �>� �)� �D ��X ��  �u� �`� �+� ��Y �:� ���  �g�  �b' ��  ��� �� �N0 �y� �d�  �o� �Z� � �@� �� �Vz �Q� �|t �GY ��I �7 �( �L �� �� �� ��� ���	 ��# ��� �[� �֥ �!a ��? ��� �{ �-X �� �� �>� �y� �t� �p	 �
� �� ��H �[� ��~ �A� �l, ��	 �2� �� � �ӭ �N �)� ��� � �j2 ��w � X �ˆ �� �!� �|� �� �b# 魀 �X1 �� �n� �I� � ��* �� 鵰 �P ��� �6� �q� ��� �g� �2� ���
 �X �#�  �>9 �		 鄊 �o@	 銢 �es �� �� �v�
 �� �\�  ��V ��  �� � ��� �>E	 �� ��/ 鏢 �j� �� �=
 �� 閗 鱥 � 	 駤 �r� �� ��@ � �� �Y� �� �O� �� �	 �d �;� �=
 ��O 鬫  ��� �2� �� �h� 铐 �^� �)6 �$� � ��� �� �s � ��� �� ��	 �$ �� �͊ ��
 ��� ��	 �)� ��E ��	 ��* �5�  ��� �[ �6- �6 �L8 闫 �r� �M�  �H� ��e �n� �yt ��� ��  ��� ��< ���	 �;H �F� �a� ��� �'8 �	 �� �hT �m �,q �Y� ��� �_� �m �u� � �� �B �AG �l� 釉 �҆ 齀 �8) �� ��� ��s	 锒 ��� �
� � ��� �� �f �a� �A	 �'9 �� ��� �ؼ ��� �� ��@ �D) �� �*� �E� �4F �+ �f� ��� �� �g�
 �� ��  �( �2 �~� 驲 �Ĭ  鯧 �7 �E�	 �о �� �� 鱲  �� �� �� �� �x� �S ��  �� ��t �o� �� ��� �L
 �� �& �a�  ��
 �� �rL �=o 騪 �R �.7 �i& � �$ �� �� ��� �\ �g �� �,� �f ��  �́ �� ��C ��d �i� �� �/� �� �5� � �� ��� �QG � �ǥ �bI �3 ��� �@ �N� ��v �$� �Z ��N ��| 頥 黊 閆 ��4 �� �� �� �M� ��j ���  �>� �� � �o �jL �5B �@�	 �{� 醱 道 �, ��v �r �� ��J
 �  ��7 �)� �TQ ��  ��� �� ��	 �� ��o �� ��/
 �W� ��{ �?	 �M ��1 ��� ��~ �C �o�	 ��j ���  �P  �� �v� 鱹
 ��  ��� �"�	 �5 �h� ��o �C �Ɏ 锤  �b �Z�
 �� ��& ��� �� �� �<% �S �� 靹 ��r ��} �>� �I� �T ��m ��! ��x �`� �Z�	 �F �!�  �� ��F	 �r� � ��a ��e �A 鉌 � �OY 銈 � 週  � �6� �!6 ��P ��� � �� � �� ��  ��� �� �O< ��  �� �  ��� �6� �\ �|x ��  �� ��&
 �H�  �#& �.�
 �y ��r �?� �: �l �p� �;� �v� �j ��/ 釒 �b7 �ݦ  �� � �� 鉓 �>	 ��� �*B �� �p� �� �v' �a
 �l� �- ���  ��# �hM �cy �n� �	w ��& �/� ��g �i	 �� �k� ��? �!G
 �h �'v ��\ �}@ ��� �F
 �nH
 �� �� �� �$ �� �h 雌 �� �u �k �'?	 �B
 靐
 � �c� ��j �y� �Ty ��	 �z� �u� �0� �kq �� �a� �L�
 � �� ��� �� ��
 �\	 �� �% ��	
 �:T �q ��) �E
 ��5 �v �\�	 �7� �r\ �� �, �c� �^� ��c ��
 �� �z
 �� �p�  ��O � �i �� ���  �,@ �M � �� �N� �	 �$a	 � �B> �} �0� �k� �fG ��7 ��� �7 �BB ��
 鈥
 鳺 �� �� ��" �� ��I �� �`� �k� ��  �a �lo ��# �2�
 �ݴ �� �s� �^�  �y� �d� �l ��q �e� � � �K-	 �V� �� 鬹 ��H 鲱  ��T ��G �( ��
 �Y� �4@ ��
 �| ��� ��( �q �Vd � �L" �= �i ��  ��� �S �nv �i ��� �?z � ��� �� �۟ �fQ �� �= 駑	 �� �m �8� �h �Ρ �	� �� �� �*� �u� � � �K	
 �v� �� �|� �$ ��P �͡
 �H� �� �) �G �^ �? �Z	 �e �� �@ ��	 �q� �Ԓ ��� ��@ �]�  �Ȇ ���	 �� ��} �$�	 ��� �J  ��� ��
 �k�  �6� �� ��� �[ �3 �_ �K �s� �� �	� �t� �y �	 �ը
 �P� �� ���  ���
 鬷 釖 �� ���  ���  �K ��e �y �d�  ��� �
� 鵹 �� �K� � �1�  � �G�
 �R�	 ��
 �H_ ��� �$ ��2 � �7
 ��  �%� � G �=	 �F �ad �\� � �B� �}D
 �ȸ �-; �~8 鹇 �l; �x �*�
 �= ��� �+ �VN
 �q�
 鬪 釣 ��* �m� ��n �3� �^4 �iy ��� �� �
� ��*	 ��� �� �Fe �1�	 �,� �� �"` ��  �c �  ��� �Y� ��� �6 �j:
 镰 �P� ��� �z 镐 ��l �� ��� �* �x� �� �>� �� ��
 �o� �0
 �� ���	 ���
 � �n �� �
 �r� �-� �(: �SY �~�	 �� ��1 �/_	 ���	 ��	 �@� �+ 鶶  ��
 ��` �w{ 邼 �J �7 ���  �.� �� �t 鯷
 �*� �u� ��$ ��� �� ��| � ��) �
 �m� �� �� 鞍 �i� �d�  �� �*� 酋 ��� 鋆
 �ֶ ��M �\� �� ��� ��  �H�
 �N�	 �ޚ ��  �4� �� �Z� �e �� 雀 閭 ��k ��  �7� �� �m� �h�  ��� �� ��� �? �~ �Z� 饊 �� ��� �6h ��	 ��� �G �"� � �8� �3& ��7 ��� � �� �j� �u�	 �� �� �f� �1� � �W! �
 �-�
 �� 鳲 �~� �9� �� ��� �Z� ��\ ��v �+~	 �� ��E ��m �� �1 ��� �(� �S� �n� 陈 ��� ��
 �Zi �� �0� �f �� ��� �� �* �h �md ��� �8 �N#
 � �D� 鯇 ��� �F �� �{� �� �A �� �7� ��� 靚 ��
 �3 鞁 �i�
 鄻 ��� �Ju �7 �X �� �V� �a� �,� � �b�  �m� 阼	 �� � 	 鹹 �� �U7 �j& �E�	 ��" �+� �v
 �1� � �G" �2� �` �� ��  �^�	 �ɷ �� �� ��$
 �D �� �e �V 
 ��  �� �' 
 �U � �(- �C� � �)�  �I �/� �: �5� �6 ��( �n �a
 �\. �� �C �� �� ��	 �!� �i� �$g �o� ��� �e� � � ��  �� �!/ �� �[ � �
 �H	 ��� 鞨 �	 �d� �b �j
 ��� � �k0 ��  ��� ���  ��� � ��� ��� �" �^�  ��� �t� �?& �*
 �E�
 �� ��3 �! �A�
 ���
 �7� �� �mH	 �hY �s �� ���	 ��z	 � � �%� ��h 鋦 �� ��� �� �� �� �� ���
 ��) �� �i� ��, �/� 銞 �%O ���  �� �V� �ag �L` ��� �b� �& �H�	 �sj �� ��� �  �?d �zt ��:
 � � �+� �Ft ��J ��� �g�
 �B �̈́ �J4 �C� �� �� ��� �� �J� �U� ��0	 ��� �� �Q� �l8 �Ƕ �"�  �` ��N �ý �>� ���	 ��  ��
 �6 ��� �@ �;o �&� �� ��� ��� ��  �-D �� �s� �.� �� ���  ��$ �� ��� �P �{/ �fQ �q �% ��� �"� �� ��+ � �� �	 �� ��� �% ��w �@6
 ��� �6 �1 �� �� �j �-�	 �H� ��	 �nZ �s �D� �o% �� ��� �7 �K� �v� �	 �|� ��. �"� �
 �X� �Ө �� �Y� �Ԩ ���  銆 ��	 �� ��  �& �a? � �e ��+ �� �([ �S� � ��� ��h � �� �� � �+� ��� �1� �� 闭	 ��  �� 鈦 �c �^� �
 �DZ ��  �e�	 ��� �0 ��# �� ���	 錂 ��	 �­ �� �(� �S�
 �N �ɢ �$� �/. �Z� ��� � �+ ���
 ��V �< �Wn �� �}� �Xe �� �s �	W �4�  ��� �z� ��� � � �� ��<	 �Q,
 � �' �2� �-� �H ��y ���	 �I�  ��z � �	 �� ��$ � 馽 �A� �۾	 �� �j 魶	 �� ��, �� 鉔 �� �? ��� �! �p� �k�  �6 �� 鼓 �G�  �R� � �X� �3 鎇  �)�	 � �� ��� �� �@
 �g �� �A: ��d �� �/ 魖	 �8� �S  �e � 鄩 韕 �� 鵟 �� �< �-
 ��,
 � �Ƕ ���  �� �(i ��y �.Q �iN �df �?` �Z� �E�	 ��v �[ �^ �As	 ��' �W� ��p	 �� �� ��� 龞 �� � 韥 �*� �E ��* �+) � ��� �, �g�	 ��  齻 � �� � ��� �t� ��� �e �5l � �/ ��. ��� �� �g� �v �Mr �s �3� ��� �z �� �V	 �� � �`f 雀 �v\ �!� �|� �	 �r� �ݷ �� 郓 ��Y � ��  ��x �*� �կ ���
 �[� 鶻 �! ��� 駱 �£ �F � �� �~ �� ��. ��$ �*� 饌 �� �{�  �f" �. 鼴 �� �� ��U ��\ �s� �N*
 ��� �$5 ��  ��� ��� � �� �FZ �!Y �Y �7P � �=*
 騾 �Y �Y ��X �� �� �:� �e� 逷 ��X �F� �] �L� �W/ �2� �� �H� ��� ��� �9� �D� �/J ��A ��T	 �@� �kd �� 遭  ��� �� �& �#
 �g 鳓 ��A �9u �h �� 骪 �P �� ��\ �6 ��P �@X �� �l �]� �X �#* �P �T	 �ċ ��
 �Z~ �eo	 �`� ��z ��W �W ��  �- ��h ��� �x: ��  �>�  �Y# �T� �O� ��( ��� �p �+�
 �v�	 ��N �|
 ��� �, ��	 �x �c
 �� �)� ��y	 ��i �Z� ��z �s
 髏 � �q� �, �G�	 �� ���	 �(�	 �7 �^� �� �� �_� �ھ �e�
 �� �[~ �f� � �, �w� ��� �-� �(� �" 龠  ��4
 �4�	 �� 麟 �՟ �{ �˒ �F �# �� �G4 � �H ��R �Cb �� �I� ��A ��^ � ��N �@z �k�
 �h �� �l*
 ��
 �� �] � �� �ާ �� �d 	 ��� �� �� �p� �N 醕  �!� �f 鷻 � �} �x� �S�  �@ �� �x	 �/� ��\ ���  �� �{� �6� �Q� 鬋 � �B� �� �X	 �� ��= ��} �dP ��	 �: �u� � | �� �V� �w) ��7
 �'� �y �� �h& �� ��u �9�  �� �_� �h �Ň �`y �[� �W �< �I �7� 钅	 �݇ �ȱ �Ê �0* �F ��� �3 �� �� ��$
 �;� � �� ��H �w� �2Q �� �~ ��	 �� �� �Dz �?� �� �$
 �Р �;� �v& �Ѩ �o ��] �b� �}�	 ��� 郟 �~� �) �4&
 ��� �Z� �EZ � ^ �� �G ��F �|< �'y
 �z 鍆 �� �� �NG	 �X ��  �� �� �� � M �1 ��( �� �� ��  �r� ��� �8a �� �>T �i| �DQ	 �?� �jH �E� �` ��8 �� ��P �\( �7� �z	 ��� �%~ �� �� �)�  �$� �� �*u �uP	 � � ��  �) �q� 鬺 ��	 �"� �=� �xu �: 铻 陻 �b �] ��� ��  � �  ��� �� ��� �\�  �%( �bu	 � �M �O �nq �� �t� �9( �*� �+
 ��� ��� �& �Qf ��  ��� �R� � � �� �& �){ �t �o)
 �:� �e� �� 馺 �� ��  �� �GV ��	 齓 �8� �cN 龫 �Y� �� �| �z�  �e�  ��� � �&� �Ai �B ��� ��c �M� �x^ �� �*
 �� ��# �� �
 �E� �� �K� ��	 �	 �|` �d �b� �g �� �C 龈 �i  �u �� �JU ��
 ���	 �{� �� �� � �� �� ��O �8� �� �>� ��	 �r ��� �*� �e� �� ��� �{ �M ��X
 �g� �P 魡 ��� �C �� ��� �X ��  �*q	 �� ��% ��� ���	 ��	 �� �W� �b�  �M� �(W �5 �N 鹝
 �t� �O�	 �_ �E� � �;� �v�	 鱹 �l� �G� ��� �ݶ �W �
 �nw �i �� �O� ���	 �Y �� ��  �� ��Q �lw	 �׉ �,% �]� �� �b �.� ��[ ��	 �o- �j�
 �5� ��n 髰 ��� �O �l� �w�	 ��� �]� �	 鳦	 �p �	� �ġ	 �Ol �:H �	% �T �KM �� �a� �� ��  �R� ��� �� �g	 ��� ��� �$�  �N �*� �}$ �J �;� �2 �!y  �z �7Q �@ �M� ��� ��? �7 �� � �F �je 酡 ��1 �{� �a ��� �lt � �� ���  �G�	 �	 ��_ ��� 餳 ��� 銵 �U�	 ��� 黈 �+ ��	 �I �4 �b� ��3 �� �4 鷱	 ��� ��4 �, �q �% �� �k �~  顪  �� ��j �? �}� �Ȱ �s�
 ��� 驊 �4� �O�	 �� ��� ��m �W ��� ��  �|0
 �g� �L �mP �H�  �I ��� �2	 ��� 鿂 �*� �Œ �. �`� 鶤 �� 錯 �� �� �}d �h� �S� �.� ��n �4y ��	 �zg �%r �@�
 ��	 �� �q ��� ��
 颦 �̓ �X �� ��� ��	 �T� �q ���	 �e� �`� �� ��� ��"	 �� ��O �2�
 �H 醯	 �s	 ���  �	� � �'
 �ZP �� �0 ��  �� 鱰 �� �� 鲭 �� �	 ��t �� �s �Dw �_X ��&
 �� �� 鋓 ��� �Q) �� �� ��& ��h �ؤ �C� ��  �I� ��� ��7 ��(
 ��' 逜 ��"	 �&�  �AJ � �g� �� ��� �8� �3w ��v �	s �4  ��

 ��( �s �P)
 �K� �Vs �a� �� �E � �Ͱ �x�  �3 �# 鉲 �l �Y �j� � �`r �{� �d 鱈  �<� ��� �b� �=� �8� ��	 �P ��t ��2 ��  �* �5� ��� �K}  �� �qr 錫 �'� ��� �=(	 �h� 郉 �� 陜 �d� �/�  �Z� �Ś �  �;� ��# �Q  �|� 鷃 �RH �mr �g �* ��e �� �tI �� �ʦ ��� �4 �� ��E �: �� �7�
 ��
 �M� ��� �w 鎛 �ɸ  锔 �� ��� 鵹 �O �� �� ��
 �1
 �G� �B 
 �� ��� �� �� �Y	 鴏  �a �� �E� �P� �� ��� � ��: � �"� �� �(� ��& ���  �Y� �h � �j�	 ���  � � �K+ �h �� �ܼ ��� ��0 �m� ��� �C� �� �Y�	 �4\ ��� �� �T �0� �� ��� ��} �<� 闣 �� 鍐 鈴 �" �N� ��  ��� �' �:  �� �0� �K ��] �1� �\�
 闏 颂  ���	 ��s �c� �ހ ��� �$� �� �:�	 �Ex �� �
 �� � �� ��� �� 齾 � �S �n� �� �4z ��x �J� ��� �� 雧 � �� �� �7a 鲬 �m� ��( �cC 龚  �y� �d�	 ��Z � �U
 �`N �˂ �ֳ �A� �{  �G� ��  ��� 鈎 �] �~N � �: � �c �%� ��� �R ��� �� �,� �G� �z ��� 騬 �� �~ ���  锨 �_� 隼 ��p �@H �;� �k � �<�  闡 � �]. �xh �k � �YM �� �� �n �5� 鰹 ��) ��� �A> �L� �W> �� �5 �H= �C�  �N� �> �m ��� �
� �E� �� ��
 ��� �q� 鼃 �K �b� ��7 �8� �� 鞖 �	� �$y �� �j� �5� �m �[� � �C �< �gI �r� �}� � �S� ��@ �9! ��  �| �ڋ �u �� ��t �� �q� �h �w� � �-� ��	 �� �� �9� ��$ ��� �z� 饉  ��I ��n �g �� ��� � �2� �� 阰	 �� �.� ��` 鴏 鏢  �
 �u�  �� �� �: �aK �� �7  �bI �M� �x* �!
 �{ �O �d�  �o� �I 酑 ��
 �� �f� 遥 �|�  �� �rd �� �R �	 �>� �9� �D� �n �T �d �`� �{ �" �� ��� �� ��� �=V ��	 � ��  �Y �4c �/P �z� �%� �p? �^�	 ��
 �qX �L ��� �
 ��- �H�	 郁 �
 �	� ��  �� 骤 �� �@�	 �� �&� �� ��� �= ��� �}5 ��� ��x � �H �k	 �} �j!
 鵍 �`� ��m �V{ ��/ �!
 �72 �� �=�	 �X� �Ә �U �c �w �? �w �� �0� �{� �m 遫 �7 �� ��	 ��	 ��P �Ý �N� �i� ��	 �/� ��� �N	 �Pt ��	 �v�	 ��j 錬 ���	 ��
 ��{  �H� �Ӭ �.�
 ��� �4� �� �ZI � �� ��O � �1x �|� 鷎 � �] ��� �s � �I� 鴮 �� �
� �Un	 � � �K �f� �
 �,� �} �
 �=q  �xS �p �~� ��	 ��L ��2 �P �� �� ��@ �� �62 ���  ��Z ��� �N �hf �� �N� �yC �! �B �2 �UT �, ��� �v� ��� �ܼ �a �J �-� 騱  �� �� �Y�  �� ��- �ZP �5�	 逦 �kW 醏 ��Y �<	 �| �� ��  �ؿ ��R �7 �� �4� �_� �Z� �E� � �	 髫 �vE �� ��	 �'j �"� ��H �8� �>A �� ��
 ��� �k 麽  �b ��� �{� �f �q� �L� ��O �b� �� �/ �#� ���  �� � �9 �� ��~ ��Y �$ �v� ��P ��� 釭 �� �=� �� �ӣ �΢
 ��S �T� �?� �Z� �� � ) �k�  �v� �!z �T �'M 邯 �- 騊 �S� 鎒  �E � ��  �J� �5� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ���������o��h +������_^[���   ;�������]������������������������U����   SVW��@����0   ���������GY��hP+�����_^[���   ;�讓����]������������������������U����   SVW��@����0   ���������y��h�+� ����_^[���   ;��N�����]������������������������U����   SVW��@����0   ������j � ��U��_^[���   ;��������]�������������������U����   SVW��@����0   ������j �����T��_^[���   ;�詒����]�������������������U����   SVW��@����0   ������j ����zT��_^[���   ;��Y�����]�������������������U����   SVW��@����0   ������j ����*T��_^[���   ;��	�����]�������������������U����   SVW��@����0   ������j �����S��_^[���   ;�蹑����]�������������������U����   SVW��4����3   ������3���;���_^[��]��������������������U����   SVW��4����3   ������3���;���_^[��]��������������������U����   SVW��@����0   ������j����U�����裇��h�+�|����_^[���   ;��Ґ����]����������������������������U����   SVW��@����0   ��������S��h@,�@|����_^[���   ;��n�����]������������������������U����   SVW��@����0   ������j ���谁��_^[���   ;�������]�������������������U���葁��h�,�{����]���������������������U�����j��h�,�{{����]���������������������U�����U��h�,�K{����]���������������������U�����u��h�,�{����]���������������������U��j ����EQ��]����������������U��j ����%Q��]����������������U��j ����Q��]����������������U��j �����P��]����������������U��Q3��E���]����U��Q3��E���]����U�칍��N|��]������������������U��Q3��E���]����U�����Yi��h-�z����]���������������������U�����S��h0-��y����]���������������������U�����Mt��hP-�y����]���������������������U��j �����O��]����������������U��j �����O��]����������������U��j ����O��]����������������U��j ����O��]����������������U��j ����eO��]����������������U��j ����EO��]����������������U��j ����%O��]����������������U��j ����O��]����������������U��j �����N��]����������������U��hp-�ux����]���������������U��Q3��E���]����U��j ����g��h�-�9x����]�������������������U��Q3��E���]����U��Q3��E���]����U��Q3��E���]����U�����g��h�-��w����]���������������������U�����rQ��h�-�w����]���������������������U�����r��h�-�{w����]���������������������U��Q3��E���]����U��Q3��E���]����U�����if��h.�+w����]���������������������U������P��h0.��v����]���������������������U�����]q��hP.��v����]���������������������U��Q3��E���]����U��Q3��E���]����U�����e��hp.�{v����]���������������������U�����P��h�.�Kv����]���������������������U�����p��h�.�v����]���������������������U��Q3��E���]����U��Q3��E���]����U��Q3��E���]����U������d��h�.�u����]���������������������U�����RO��h�.�u����]���������������������U������o��h/�[u����]���������������������U��Q3��E���]����U��h0/�%u����]���������������U��d���z��hP/��t����]���������������������U��Q3��E���]����U������c��hp/�t����]���������������������U�����RN��h�/�t����]���������������������U������n��h�/�[t����]���������������������U��j � ��J��]����������������U��j �|��eJ��]����������������U��j ����EJ��]����������������U��j ����%J��]����������������U��Q3��E���]����U��Q3��E���]����U������b��h�/�s����]���������������������U�����"M��h�/�[s����]���������������������U�����m��h0�+s����]���������������������U��j ����UI��]����������������U��j ����5I��]����������������U��j ����I��]����������������U��j �����H��]����������������U��j �����H��]����������������U��j ����H��]����������������U��j ����H��]����������������U��j ����uH��]����������������U��j ����UH��]����������������U��j ����5H��]����������������U��j ����H��]����������������U��j �����G��]����������������U��j �����G��]����������������U��j ����G��]����������������U��j ����G��]����������������U��j ����uG��]����������������U��j ����UG��]����������������U��j ����5G��]����������������U��j ����G��]����������������U��j �����F��]����������������U��j �����F��]����������������U��j ����F��]����������������U��j ����F��]����������������U��j ����uF��]����������������U��j ����UF��]����������������U��Q3��E���]����U��Q3��E���]����U������^��h00�o����]���������������������U�����RI��hP0�o����]���������������������U������i��hp0�[o����]���������������������U��j �P��E��]����������������U��j �T��eE��]����������������U��j �X��EE��]����������������U��j �\��%E��]����������������U��j �d��E��]����������������U��j �`���D��]����������������U��j �����D��]����������������U��j ����D��]����������������U��j ����D��]����������������U��j ����eD��]����������������U��j �h��ED��]����������������U��j �l��%D��]����������������U��Q3��E���]����U��Q3��E���]����U������\��h�0�m����]���������������������U�����"G��h�0�[m����]���������������������U�����g��h�0�+m����]���������������������U��j ����UC��]����������������U��j ����5C��]����������������U��j ����C��]����������������U��j �����B��]����������������U��Q3��E���]����U��Q3��E���]����U����   SVW��@����0   ������E���Ex��M�U;��{����EE�E��_^[���   ;��`�����]� �����������������������U����   SVW��@����0   ������_^[��]������������U����   SVW��<����1   ������E��<�����<���t����~B����u3��3�_^[���   ;������]�����������������������U����   SVW��@����0   �������n�����u3���   _^[���   ;��c����]�����������������������������U����   SVW��@����0   ������E;Et��EPj �MQ�k����_^[���   ;���~����]�����������������������������������U����   SVW��4����3   �������E�    �} u� �}�w�EP�!Y�����E��}� u�O���E�_^[���   ;��s~����]�����������������������������U����   SVW��4����3   �������E�    �} u�&�}���w�E��P�X�����E��}� u�O���E�_^[���   ;���}����]���������������������������������������U����   SVW��4����3   �������E�    �} u�$�}UUUwkE0P�X�����E��}� u�~N���E�_^[���   ;��_}����]�����������������������������������������U����   SVW��@����0   ������} t#��j �E��M���;���|���EP蔇����_^[���   ;���|����]��������������������������������������U����   SVW��@����0   ������} t#��j �E��M���;��x|���EP������_^[���   ;��\|����]��������������������������������������U����   SVW��@����0   ������} tj �M�f>���EP衆����_^[���   ;���{����]�����������������������������������U����   SVW��@����0   ������} u�EP�MQhq��d����_^[���   ;��z{����]��������������������U����   SVW��@����0   ������} u�EP�MQhq�bd����_^[���   ;��{����]��������������������U����   SVW��@����0   ������} u�EP�MQhq�d����_^[���   ;��z����]��������������������U����   SVW��@����0   ������} u�EP�MQhq�c����_^[���   ;��Zz����]��������������������U����   SVW��@����0   ������E;EtE�EP�MQ�UR�}�����EP�MQ�UR��|�����E;Es�EP�MQhPq�c����_^[���   ;���y����]����������������������������������U����   SVW��@����0   ������E;EtE�EP�MQ�UR�ǌ�����EP�MQ�UR賌�����E;Es�EP�MQhPq�pb����_^[���   ;��(y����]����������������������������������U����   SVW��@����0   ������E;EtE�EP�MQ�UR�X�����EP�MQ�UR�X�����E;Es�EP�MQhPq��a����_^[���   ;��x����]����������������������������������U����   SVW��4����3   ������EP��;���Q�9o�������P�MQ�UR�EP�MQ�F����_^[���   ;��x����]������������������������������U����   SVW��4����3   ������EP��;���Q��e�������P�MQ�UR�EP�MQ�I����_^[���   ;��w����]������������������������������U����   SVW��4����3   ������EP��;���Q�3Q�������P�MQ�UR�EP�MQ��T����_^[���   ;��w����]������������������������������U����   SVW��4����3   ������EP�MQ��g������;�����;���R�EP�MQ�UR�nl����_^[���   ;��v����]�����������������������������U����   SVW��@����0   �������	�E��0�E�E;Et�EP�M�?D����_^[���   ;��v����]������������������������������U����   SVW��4����3   ������EP�96�����E��}��u2���
�E�M���_^[���   ;��u����]��������������������������U����   SVW��<����1   ������EP�MQ�s6�������tǅ<���   �
ǅ<���    ��<���_^[���   ;��#u����]�����������������������������U����   SVW��4����3   ������E�M���ER��P�t�腈��XZ_^[��]ÍI    |�����   ��_Cat �����������������������������������U����   SVW��4����3   ������E�M���ER��P�������XZ_^[��]ÍI    ������   �_Cat �����������������������������������U����   SVW��4����3   ������E�M���ER��P�t�腇��XZ_^[��]ÍI    |�����   ��_Cat �����������������������������������U����   SVW��4����3   ������E�R��P�������XZ_^[��]ÍI    ������    �_Cat ���������������������������U����   SVW��4����3   ������E�R��P�\�蝆��XZ_^[��]ÍI    d�����   p�_Cat ���������������������������U����   SVW��@����0   ������E�M��E_^[��]�����������������U���   SVWQ�� ����@   ������Y���3ŉE��M�E�P�M���G���E�P�M Q���̍UR�b�����̍EP�b���wG���� ������M��i���M��i�������R��P���荅��XZ_^[�M�3���U����   ;��q����]� ��   ������   ��_Alval �����������������������������������������������������������������U����   SVWQ��$����7   ������Y���3ŉE��M�E�P�M���F���E�P�MQ�UR�EP��p����R��P�d�譄��XZ_^[�M�3��U�����   ;���p����]� ��   l�����   x�_Alval �������������������������������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��4����3   ������M������8����M�h����8���_^[���   ;���o����]�����������������������������������U����   SVW��<����1   ������EP�M�R�`�������tǅ<���   �
ǅ<���    ��<���_^[���   ;��qo����]���������������������������U����   SVW��4����3   ������EP�MQ�|W������;�����;���R�EP�MQ�UR�EP��/����_^[���   ;���n����]�����������������������������������������U��j�h��d�    PQ���   SVW��$����3   �����󫡀�3�P�E�d�    �e�ht  h�q�EP�MQ�3����hu  h�q�EP�Mq�����E�E��E�    ��E��0�E�M��0�M�E;Et�EP�MQ�M�,~�����0�	�E��0�E�E�;Et�E�P�M�<����j j �\f���W���E�������E������E�M�d�    Y_^[���   ;��m����]���������������������������������������������������������������������������������U����   SVW��4����3   ������EP�MQ�L^������;�����;���R�EP� w����P�MQ�UR�EP�MQ�w����_^[���   ;���l����]��������������������������������������������U��j�h�d�    PQ���   SVW��$����3   �����󫡀�3�P�E�d�    �e�h�  h�q�EP�MQ�:����h�  h�q�EP�Mo�����E�E��E�    ��E��0�E�M��0�M�E;Et�EP�MQ�M�!U�����0�	�E��0�E�E�;Et�E�P�M�:����j j �\d���W���E�������E������E�M�d�    Y_^[���   ;��k����]���������������������������������������������������������������������������������U����   SVW������9   ������E$P�M Q�O����P���̍UR�[���7x����P���̍EP�[��� x����P��T����P�M Q�:f������� ����M��b���M��b���� ���_^[���   ;���j����]���������������������������������������������U����   SVW��@����0   ������EP�MQ�4N����P�UR�'N����P�EP�N����P�P����P�MQ�~e����� _^[���   ;��#j����]���������������������������������������������U����   SVW��@����0   ������3�_^[��]����������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVWQ��4����3   ������Y�M��EP�~����P�MQ�U�R�|\����_^[���   ;���h����]� ��������������������������U����   SVWQ��$����7   ������Y�M��EPj��L������,�����,��� t$�MQ��}������,���� ���,�����$����
ǅ$���    _^[���   ;��Uh����]� ��������������������������������������������U����   SVW��@����0   ������EP�i}����P�MQ�M�"K��_^[���   ;���g����]����������������������U����   SVWQ��4����3   ������Y�M��EP�i1����P�MQ�U�R�+����_^[���   ;��sg����]� ��������������������������U����   SVWQ��$����7   ������Y�M��EPj�xK������,�����,��� t*�MQ��0������@��,�����A��,�����$����
ǅ$���    _^[���   ;���f����]� ��������������������������������������U����   SVW��@����0   ������EP�N0����P�MQ�M�cL��_^[���   ;��\f����]����������������������U����   SVWQ��4����3   ������Y�M��EP�IR����P�MQ�U�R�F����_^[���   ;���e����]� ��������������������������U����   SVW��@����0   ������EP��Q����P�MQ�M��=��_^[���   ;��e����]����������������������U����   SVWQ��4����3   ������Y�M��EP�-����P�MQ�U�R�*q����_^[���   ;��#e����]� ��������������������������U����   SVWQ��$����7   ������Y�M��EPj0�(I������,�����,��� t)�MQ�)-�����   ����,���󥋕,�����$����
ǅ$���    _^[���   ;��d����]� ���������������������������������������U����   SVW��@����0   ������EP�,����P�MQ�M�(b��_^[���   ;��d����]����������������������U����   SVWQ��4����3   ������Y�M��EP�M�Q��:����_^[���   ;��c����]� �����������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVW��@����0   ������EP�M�]\��_^[���   ;��c����]�������������������U����   SVWQ��4����3   ������Y�M��EP�M�Q�I=����_^[���   ;���b����]� �����������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVW��@����0   ������EP�M�P��_^[���   ;��)b����]�������������������U����   SVWQ��4����3   ������Y�M��EP�M�Q�5B����_^[���   ;���a����]� �����������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVW��@����0   ������EP�M��M��_^[���   ;��9a����]�������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E_^[��]�������������������������U���   SVW�������H   �����󫡀�3ŉE�j �M��v1�����E� ��-���E܋E�P�M��T���EЃ}� t�|�}� t�E�E��n�EP�M�Q�H�������u#hDq�������6��hPP������P�W���6�E�EЋE���E�EċEċ��MċB��;��_���E�P�Jb�����EЉ������M�� \��������R��P�p	�r��XZ_^[�M�3��C����   ;���^����]�   x	����   �	����   �	_Psave _Lock �����������������������������������������������������������������������������������U���   SVW�������H   �����󫡀�3ŉE�j �M���/�����E蹨���+���E܋E�P�M�-S���EЃ}� t�|�}� t�E�E��n�EP�M�Q�W�������u#hDq��������4��hPP������P�V���6�E�EЋE���E�EċEċ��MċB��;��u]���E�P�`�����EЉ������M��`Z��������R��P�	��p��XZ_^[�M�3��nA����   ;��']����]�   	����   7	����   0	_Psave _Lock �����������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��U���M���E�_^[���   ;��c\����]�����������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@   �M��mX���E�_^[���   ;���[����]����������������������������U����   SVWQ��4����3   ������Y�M��M��_���E�_^[���   ;��[����]�������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���I���E�_^[���   ;��1[����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��D^���E�_^[���   ;���Z����]�������������������������������U����   SVWQ��4����3   ������Y�M��M���2���M��E���E�_^[���   ;��mZ����]� ��������������������U����   SVWQ��4����3   ������Y�M��M���V���EP�M���X���E��M�H�E�_^[���   ;�� Z����]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M��$���E�_^[���   ;��Y����]� ��������������������U����   SVWQ��4����3   ������Y�M��M��YS���E��@    �E��@    �E�_^[���   ;��1Y����]���������������������������U����   SVWQ��4����3   ������Y�M��M��f���M��)���E�_^[���   ;���X����]� ��������������������U����   SVWQ��4����3   ������Y�M��EP�M��V'���E��M�Q�P�E�_^[���   ;��eX����]� ����������������������������U����   SVWQ��4����3   ������Y�M��M��H#���E��M�H�EP�M��V���E�_^[���   ;���W����]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M��uK���E�_^[���   ;��W����]� ��������������������U����   SVWQ��4����3   ������Y�M��M��IQ���E��@    �E��@    �E��@    �E�_^[���   ;��W����]���������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���9���E�_^[���   ;��V����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��!a���E�_^[���   ;��UV����]�������������������������������U����   SVWQ��4����3   ������Y�M��M���0���E�_^[���   ;���U����]�������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���<���E�_^[���   ;��U����]� ������������������������U����   SVWQ��4����3   ������Y�M��M���+���E�_^[���   ;��5U����]�������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@ �E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��E��     3��M�f�A�E�_^[��]������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��M��U���E�� Lej �EP�M���"���E�_^[���   ;���R����]� �������������������������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �} t�E�� �e�M���p�S����,���j j �E���P�M��~:���E���Q�E���e�E���Q��p�E���A�M��T�j �M����;���EP�M��Q�UR�M�����&����uj j�E���U�Q����c���E�_^[���   ;���Q����]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��f!���E�� �d�E�_^[���   ;��LQ����]����������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �} t�E�� �d�M���������,����E���Q�E���d�E���Q���E���A�M��T��E��@    �@    �EP�MQ�U���M�H�>���E�_^[���   ;��|P����]� ���������������������������������������������������U����   SVWQ��$����7   ������Y�M��E��  ejh@m�I��Pj�d������,�����,��� t��,����[����$����
ǅ$���    �E���$����H4�M��6���E�_^[���   ;��O����]���������������������������������������U����   SVWQ��(����6   ������Y�M���/���P�M��S��P�M����j j �M���$���EP�MN����P�M�����E�_^[���   ;��O����]� �������������������������������������������U����   SVWQ������9   ������Y�M���/���P��#���Q�M�S�����wR��P�M����j j �M��J$���@aPj �MQ�M���M���E�_^[���   ;��gN����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M���/����X��P�M��e��j j �M��#���EP�MQ�M��F���E�_^[���   ;���M����]� �����������������������������������U����   SVWQ��(����6   ������Y�M���/����.X��P�M�����j j �M��#���EP�M�����E�_^[���   ;��AM����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M���/����W��P�M��E��j j �M��"���E�_^[���   ;��L����]�����������������������U����   SVWQ��4����3   ������Y�M��EP�M��E&���E�� �h�EP�M�����E�_^[���   ;��LL����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��t:���E�� �b�EP�M��=���E�_^[���   ;���K����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E��     �@    �E��M�H�U�P�E��M�H�E�_^[��]� �������������������������U����   SVWQ��4����3   ������Y�M��E��M��U�P�E��@    �@    �E��@    �E�_^[��]� ������������������������U��j�h@�d�    PQ���   SVWQ�������?   ������Y���3�P�E�d�    �e��M荅���P������Q�M�< �����D��P�M��s$���M�W��P�M��E������t]�E�    �E�HQ��T�M��!����T�M�!.���M�����U�B��M��!��j j �iB���J	��E�������E������E�M�d�    Y_^[��  ;���I����]� ���������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M���/�������P�M��X#���E�_^[���   ;��)I����]�����������������������������������U����   SVWQ��4����3   ������Y�M��M��2���E�� ,`�E�_^[���   ;��H����]����������������������U����   SVWQ��4����3   ������Y�M��E��E� �E��E�@�E��E�@�E�_^[��]� ���������������������������U����   SVWQ��4����3   ������Y�M��M��3���E�� �e�E�_^[���   ;���G����]����������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��G����EPj��MQ�U�R����H�Q�҃�;��kG���E�_^[���   ;��XG����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;���F���E�_^[���   ;���F����]�������������������������U����   SVWQ��4����3   ������Y�M��E��     �E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E�� la�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��M��=���E�� Xc�E�_^[���   ;��|E����]����������������������U����   SVWQ��4����3   ������Y�M��M��+ ���E�� �c�E�_^[���   ;��E����]����������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �EP�M��&���E�_^[���   ;��D����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVWQ�� ����8   ������Y�M�j �M������M����bA���M����WA���M����P���M����P���M���$�6A���M���,�+A���} u!hTa��$������h\O��$���P�<���EP�M�Q�Y�����E�_^[���   ;��zC����]� �������������������������������������������������U����   SVWQ��,����5   ������Y�M��E��M��E����0�����0������0���H������tC�E����0�����0������0���H�����,�����,������,����B��;��B���E�_^[���   ;��B����]� ����������������������������������������������������U����   SVWQ��,����5   ������Y�M��E��M��E����0�����0������0���H������tC�E����0�����0������0���H������,�����,������,����B��;���A���E�_^[���   ;��A����]� ����������������������������������������������������U����   SVWQ������?   ������Y�M����̋EP����MQ�UR�����P�1����(P�M��2U�����������E�� 4c�E��M�H�U�P�E�_^[���   ;���@����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��&���E�� 4c�E�H�P�E��H�P�E�_^[���   ;��v@����]� �����������������������������U����   SVWQ��4����3   ������Y�M��M�����E�� �c�E�_^[���   ;��@����]����������������������U����   SVWQ��4����3   ������Y�M��EP�M��8!���E�� �a�E�_^[���   ;��?����]� �������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��� ���E�� �b�E�_^[���   ;��8?����]� �������������������������������U����   SVWQ��4����3   ������Y�M��E�� c�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E��M��E��M�H�E�_^[��]� ����������������U����   SVWQ��4����3   ������Y�M��E��M��E��M�H�E�_^[��]� ����������������U����   SVWQ��4����3   ������Y�M��M�� ���E�� �a�EP�M���Q������E�_^[���   ;���=����]� ��������������������������������U����   SVWQ��4����3   ������Y�M��EP�M���&���E�� d�E�_^[���   ;��X=����]� �������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�QR�P�M��7���E�� d�E�_^[���   ;���<����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��E�_^[��]� �������������������������U����   SVWQ��4����3   ������Y�M��E��  d�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E��M���E���U����
�P��;���;���E�_^[���   ;��;����]� ��������������������������������U����   SVWQ��4����3   ������Y�M�j�,�����M���E�_^[���   ;��N;����]������������������������U����   SVWQ��4����3   ������Y�M��E��E� �E��E�@�E��E�@�E�_^[��]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�M��cC���E�� Ha�E�_^[���   ;��x:����]� �������������������������������U����   SVWQ��(����6   ������Y�M��M�����,�����,���P�M�����E�� Ha�E�_^[���   ;���9����]� ������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��N���E�� Ha�E�_^[���   ;��9����]� �������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�����EP�M��	�)I���U��B�E�_^[���   ;��9����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��l���E��UQ����������tF�E��UQ���l(����t0�E��UQ���V(��;Et�E��UQ���?(������3���E��UQ���2����M��A�E�_^[���   ;��*8����]� �������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M������E��P�M��������E�_^[���   ;��7����]� ����������������������U����   SVWQ��4����3   ������Y�M��EP�M�����M����#���M�
���E�_^[���   ;��.7����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M������E�� Hc�E�_^[���   ;��6����]� �������������������������������U����   SVWQ������<   ������Y�M��EP������>�������Q�UR�EP�M��j��������	���E�� Hc�E�_^[���   ;��#6����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��U�P�M�H�E����M��U�P�M�H�E����M,��U0�P�M4�H�E���$�M ��U$�P�M(�H�E�_^[��]�0 ����������������������������������������U����   SVWQ��4����3   ������Y�M��E�P�D�����E��     _^[���   ;���4����]���������������������U����   SVWQ��4����3   ������Y�M��M�� 1��_^[���   ;��4����]������������������U����   SVWQ��4����3   ������Y�M��M��[��_^[���   ;��X4����]������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;��4����]������������������U����   SVWQ��4����3   ������Y�M��M��)���M��dD��_^[���   ;��3����]��������������������������U����   SVWQ��4����3   ������Y�M��M��;��_^[���   ;��X3����]������������������U����   SVWQ��4����3   ������Y�M��M��z���_^[���   ;��3����]������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;��2����]������������������U����   SVWQ��4����3   ������Y�M��M��\���M��P���_^[���   ;��`2����]��������������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��2����]������������������U����   SVWQ��4����3   ������Y�M��M���)��_^[���   ;��1����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��h1����]������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;��1����]������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;���0����]������������������U����   SVWQ��4����3   ������Y�M��E�� Le�E��xP t�M�����E��HL��t�M��_ ���M������_^[���   ;��K0����]�������������������������������������U����   SVWQ��4����3   ������Y�M��E��H��Q�E��D��e�E��H��Q��p�E��H��A�M��T��M���`�4>���M���X����_^[���   ;��/����]������������������������������������U����   SVWQ��4����3   ������Y�M��E�� �d�M����_^[���   ;��?/����]�������������������������U����   SVWQ��4����3   ������Y�M��E��H�Q�E��D��d�E��H�Q���E��H�A�M��T�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��E��  e�E��H4Q�G�����_^[���   ;��h.����]����������������������������������U����   SVWQ��4����3   ������Y�M�j j�M������M��"��_^[���   ;���-����]����������������������U����   SVWQ��4����3   ������Y�M��E�� �h�M��U��_^[���   ;��-����]�������������������������U����   SVWQ��4����3   ������Y�M��E�� �b�M��"#���M�����_^[���   ;��7-����]���������������������������������U����   SVWQ��4����3   ������Y�M��M�����M�����_^[���   ;���,����]��������������������������U����   SVWQ��4����3   ������Y�M��M��,��_^[���   ;��x,����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��(,����]������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;���+��_^[���   ;���+����]����������������������������U����   SVWQ��4����3   ������Y�M��M��s��_^[���   ;��h+����]������������������U����   SVWQ��4����3   ������Y�M��E�� la_^[��]��������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;���*����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��*����]������������������U����   SVWQ��$����7   ������Y���3ŉE��M�j�M������M��o���M��4'��R��P�86	��=��XZ_^[�M�3��H�����   ;��*����]Ë�   @6	����   L6	_Lock ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E�P�-�����M���,�m+���M���$�b+���M����_���M����T���M����A+���M����6+���M��B&��_^[���   ;��*)����]������������������������������������U����   SVWQ��,����5   ������Y�M��E����0�����0������0���H������tC�E����0�����0������0���H�r�����,�����,������,����B��;��x(��_^[���   ;��h(����]��������������������������������������������������U����   SVWQ��,����5   ������Y�M��E����0�����0������0���H�������tC�E����0�����0������0���H������,�����,������,����B��;��'��_^[���   ;��'����]��������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��('����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;���&����]������������������U����   SVWQ��4����3   ������Y�M��E�� �a�M�����_^[���   ;��&����]�������������������������U����   SVWQ��4����3   ������Y�M��E�� �b�M��9���_^[���   ;��&����]�������������������������U����   SVWQ��4����3   ������Y�M��E�� c_^[��]��������������U����   SVWQ��4����3   ������Y�M��E�� �a�M��k��_^[���   ;��%����]�������������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;��(%����]������������������U����   SVWQ��4����3   ������Y�M��E��  d�E�P������_^[���   ;���$����]���������������������U����   SVWQ��4����3   ������Y�M��E��8 t#�E���U����
�P��;��n$��P�������_^[���   ;��U$����]�������������������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;���#����]������������������U����   SVWQ��4����3   ������Y�M��M��8��_^[���   ;��#����]������������������U����   SVWQ��4����3   ������Y�M��������u
�E����/���M�����_^[���   ;��B#����]����������������������������U����   SVWQ��4����3   ������Y�M��M����H����M��`���_^[���   ;���"����]�����������������������U����   SVWQ��4����3   ������Y�M��M��]���_^[���   ;��"����]������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������EP�MQ�UR�EP�
6����_^[���   ;���!����]�����������������������U����   SVW��@����0   ������EP�0�����_^[���   ;��!����]�������������������U����   SVWQ��$����7   ������Y���3ŉE��M�E�M�;u�4�E�8 t�E��R�M������j�M�������M��W����M�����E�R��P�T?	�4��XZ_^[�M�3��-�����   ;��� ����]� �   \?	����   h?	_Lock ��������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��y��_^[���   ;��X ����]������������������U����   SVWQ��0����4   ������Y�M��EP�M���	���E��M�P;Quǅ0���   �
ǅ0���    ��0���_^[���   ;�������]� ���������������������������������U����   SVWQ��0����4   ������Y�M��E�;Euǅ0���   �
ǅ0���    ��0���_^[��]� ��������������������������������U����   SVWQ��0����4   ������Y�M��M���P�M�������B������t"�M��������M����;�uǅ0���   �
ǅ0���    ��0���_^[���   ;������]� ��������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��}#���ȅ�uǅ0���   �
ǅ0���    ��0���_^[���   ;��1����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|.h,hh�   hHhh�h������hHhh�   �=/�����E��H�U��_^[���   ;������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��Q�pq��_^[��]������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��$����7   ������Y���3ŉE��M�E�8 u2j �M��I����E�8 u���������M�����M��d���E� R��P�D	�0��XZ_^[�M�3��s �����   ;��,����]Ð   D	����    D	_Lock ����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��M��|�����tD�E��x t;�M��g���������M�9Ar$�M��P������i�����M��?���p�E�;pw_jOh�fh�o��������i��t3�u#hjhpjj jPh�fj���������u�j jPh�fh ph�k������E��@_^[���   ;��+����]���������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;������]������������������U����   SVWQ��4����3   ������Y�M��M��������t/�E��x t&�M�������M��Q;Pr�M�������M��P;Qw_jHh�hh�i�Y������i��t3�u#hjhpjj jIh�hj�g�������u�j jIh�hhxjh�k������E��@_^[���   ;�������]����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;��H����]������������������U����   SVWQ��4����3   ������Y�M��M�������t�E��x t�M������M��P;Qw_jeh�hh�k�������i��t3�u#hjhpjj jfh�hj��������u�j jfh�hh lh�k�������E��H��0�U��J�E�_^[���   ;��g����]�����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�����E�_^[���   ;�������]�������������������������������U����   SVWQ��4����3   ������Y�M�j�j��EP�M��o#��P�M��~���E�_^[���   ;��t����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M���p�&���M���p���_^[���   ;��
����]��������������������U����   SVWQ��4����3   ������Y�M��M���������M����[��_^[���   ;������]��������������������+I��v����+I��8����������������U����   SVWQ��4����3   ������Y�M��M��#���E��t�E�P�)�����E�_^[���   ;��!����]� ������������������������U����   SVWQ��4����3   ������Y�M��M���p����E��t�E���pP�(�����E���p_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�$(�����E�_^[���   ;��1����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��������E��t�E���P�'�����E���_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�4'�����E�_^[���   ;��A����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��Y����E��t�E�P�������E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M��F'���E��t�E�P�C������E�_^[���   ;��a����]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P��%�����E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�t%�����E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�%�����E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�$�����E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�$$�����E�_^[���   ;��1����]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�#�����E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M��r$���E��t�E�P�D#�����E�_^[���   ;��Q����]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P��������E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�S������E�_^[���   ;��q����]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P��!�����E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�s������E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�!�����E�_^[���   ;��!����]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P� �����E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M��G����E��t�E�P�4 �����E�_^[���   ;��A����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��S����E��t�E�P�������E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�T�����E�_^[���   ;��a����]� ������������������������U����  SVWQ��@�����   ������Y���3ŉE��M�j�M�������M�����j h�e��`����*�����H������P��`���Pj j�M��������H����������`��������j hf�����������������P�M��������x���������������x��� �  j�M��'����M������h1D4ChCD4Cjjj�E�P�M���������Z�����u%ǅ����    �M������M�������������  j�M����j h�a�M��?����M��������h����E�ǅ����   ������s��"���������D� �   k� �T��U�ǅ|���    ���|�������|�����|���;E�tE�E�P�M������������j �E�P����������P�M������������v�����|���~��j hf�������|���j j ������P�M��I�����t	ƅC����ƅC��� ��C�����s��������������M�������������s������7  j ������P�M�����������P�� ����{���� ���Q��<���R�������� ������������������M��x��j��$���������$���P�M�����j������������X���P���������ǅ ���    ǅ����    ��X���������j�����������������P����������j����������������P������������������Y���������P��������
���ȅ��E  �������w����   ����������Z��������$�Z��������$�Z��������$��h��������Z��������$�Z��������$�Z��������$��H����l����Z��������$�Z��������$�Z��������$��(����1���jj�������� ����� �������������� �������������   k� ������h������l����A��p����Q��t����A��x����Q��|����A�   �� ������H������L����P��P����H��T����P��X����H��\����P�   ��������(������,����P��0����H��4����P��8����H��<����P������     ������@   ������@   j j�� ���������� �����������$���P���������������P����-���j j j �� ���P�M�[���������������������������ǅ���    �����������������+���9����}j�����P��������������j h�A  �J����j h�6  �;����j ����������]����X���������<���������������������������$����������<����'����.j hf�����������j0������P�����������������M������M������j �3�����ǅ���   �M����������R��P�\	����XZ_^[�M�3��m������  ;��&����]� �   \	����   �\	����   �\	����   �\	����   �\	<���,   �\	$���   �\	���   �\	����   �\	����   �\	����0   �\	h���   �\	H���   �\	(���   �\	c b a t $S3 $S2 triangles name info c text bf file �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M��B@��;��� ��_^[���   ;��� ����]� ����������������������������������U����   SVWQ������9   ������Y�M��E��8 tD�E�    �E��H�M��E�    ��E���E�M����M��E��M�;H}��E�P��������E��     �E��@    �E��@    �E��@    �E��@    _^[���   ;�� ����]�������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M�����P��M��B<��;��W���_^[���   ;��G�����]���������������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M�����_^[���   ;��������]���������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M�����_^[���   ;�������]���������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���   �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M��} }3��.jjj�EP�M�������u3���E��H�U�E���   _^[���   ;��x�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M��BL��;�����_^[���   ;��������]� �����������������������������U���P  SVWQ�������T   ������Y�M��} }3��t  �} 
�   �d  �E��H;M~�U��B�������	�M������������U�U�E��x uhHhhA  ������3��  �E��H��9M��  �E��H+M�U��J�E��x ��  �E��@�؃��M���y���U��B��E܉U��E��@�E�U�j jRP�_���ẺUЋE̙�������������E�;�����ud�M�;�����uY�E��@�E�U��������������M�;�����|5�U�;�����r(�E��������������E�;�����K|�M�;�����s>�   ��t.h�qhP  hHhh�h�B�����hHhhP  �����3���  �E܋M�A�U��B�E܋M�A�U��B�E��8 u8��hHhhW  �E��H��Q����B���  �у�;�������U���<��hHhhX  �E��H��Q�U��P����Q��  �Ѓ�;������M���E��8 u3��@  �E��H�U�����U��J�} ��   �E��H+M��Q�E��ȋ�+M�u��E���j jVQ����U�BP�EE�M��Q��P�������E��P�E�+E�U�j jRP�l���M�AP�U��BP��������;�E��H��Q�E�+E�U�j jRP�5���U�BP�E��H�U��P�������?�} ~%�E��P�M��QR�E��H�U����Q�u������E��H�U�����U��J��  �E��H�U�D
��M���y���U��B��E��U��E��@��������������M�;������g  �U�;������V  j j�E�P�M�Q�j���E��U��E���������������E�;�����uE�M�;�����u:�E�;E�|2�M�;M�r(�E��������������E�;�����K|�M�;�����s>�   ��t.h�qhx  hHhh�h�l�����hHhhx  ��	����3��  �E��8 u5��hHhh|  �E���P����Q���  �Ѓ�;������M���8��hHhh}  �E���P�M��R����H��  �҃�;�������M���E��8 u3��  �E��H�U�����U��J�E��M��A�E��M;H}2�E��H+M��Q�U��B�M��R�EE�M��Q��P�q������E�    �E�    �} ti�E��H;M}5�E��H�U��B��Q�U��E+B��P�M��Q�E��H��R�������E��H�U��P�M��Q�U��B�M��R��������} ��   �E��H;M}M�E��H�M��U��B�M��Q���E���E����E��M����M��E�;E}�E�Pj����������������E�    �E��H�U���E���E����E��M����M��E�;E}�E�Pj�������������ЋE��M�H�   _^[��P  ;�������]� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ������   �M��P��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��HQ�UR�M�葿��_^[���   ;�������]� ��������������������U����   SVWQ��4����3   ������Y�M��E��M;Hu�   �@�E��M;H}�E��H+MQ�UR�M��(����jj�E��M+HQ�U��BP�M�����_^[���   ;��������]� �������������������������������������U���  SVW�������F   ������hHf� ���Ph�j������������������� t�������7����������
ǅ����    j h�f��,�������������Qj h�f������y���P��,���R�� ����5���������Pj h'  �����Ph@B �:������������� �������������� �����,��������������_^[��  ;��������]����������������������������������������������������������������������U���  SVWQ�������E   ������Y�M��} 
�   ��  �} |�E��M;H}�E��8 u3���  �E��x uhHhh�  �����3��  �} �E��M;H|�M��]����   �  �E��HQ�UUR�	������E�E�+E�E��E�    �E�    �E�    �E��H�U���E���Eԃ��EԋMȃ��MȋE�;E�}��E��H��9M�"  �E��HM��U��J�} ~#�E��P�M��QR�E��H�U���P�K������E��H�U�����U��J�E��M��P;Q��   �E��M��@��y�U��B�E��E��H+M��U��J�E��H+M��U��J�E��H+M���Q�U��BP�M��ًU��B��Q�Ž������hHhh�  �E��H��Q�U��P����Q��  �Ѓ�;������M���E��8 u3��  �E��H�U�����U��J��   �E��H�U��B�D�+E��M���y���U��B�E��E��H��9M}7�EE��M��Q+���R�EE��M��Q��P�M��Q�E��Q��������E��M�;H}a��hHhh�  �E���P�M��R����H��  �҃�;������M���E��8 u3��1�E��H�U�����U��J�E��M��H�E��H+M��U��J�   _^[��  ;��X�����]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q@�B�Ѓ�;��B���E��P�M�Q����B@�H�у�;�� ���_^[���   ;�������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��B|��;�����_^[���   ;�������]� ����������������������U����   SVW��@����0   ������E;E}�E��E_^[��]����������������������������U����   SVWQ������=   ������Y���3ŉE��M�} uj�M�諽���M������M�������I�E��M܋E�;M�t7j�M��}����M�������E�M܋Q�P�E܋M�H�E�M܉�M�����R��P��t	�6���XZ_^[�M�3��������   ;��`�����]� �I    �t	����   u	����   �t	_Lock _Lock ������������������������������������������������������������������������U����   SVWQ������;   ������Y���3ŉE��M�M�����j�M��u����M����������P�E�Q�M��|����E��U�R��P��u	�&���XZ_^[�M�3��������   ;��P�����]Ð   �u	����   �u	_Alproxy �����������������������������������������������������������U����   SVWQ������;   ������Y���3ŉE��M�M��&���j�M��n����M����������P�E�Q�M��
����E��U�R��P��v	�6���XZ_^[�M�3��������   ;��`�����]Ð   �v	����   �v	_Alproxy �����������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�xs"�E�H��Q�U��R�E���P聸�����.�E��P�M���Q��/���R�M��������:����E�@    �E��M�Q�P�E��M�Q�Pj j �M����_^[���   ;��S�����]� ����������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��@    �E��@    �E��@    �} u2��W�S�M�����;Es
�M�������<�EP��/���Q�M��q����������U��B�E��M��Q�PkE0�M�A�U��B�_^[���   ;��a�����]� ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M��}u�EP�M�����EP�*�������EP�MQ�M�����EP�!�����_^[���   ;�������]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     _^[��]��������������U����   SVWQ��4����3   ������Y�M��M�謶����t�M�蠶�����M薶��;�thh�   h�hh�m��������m��t3�u&h(nhpjj h�   h�hj�*�������u�j h�   h�hh�nh�o�������_^[���   ;�������]� �������������������������������������������������������������U��j�hp�d�    PQ��  SVWQ�������C   ������Y���3ŉE�P�E�d�    �e��M�E���E؋M��m���;E�s�E�E��R�E�H��E�3Ҿ   ��;�w�8�M��>����M�Q��+M�9Aw�E�H��U�J�M���M������E��E�    �E؃�P������Q�M��������軭���E��`�e��E�E��E��E؃�P������Q�M�������茭���E��j j�M�����j j �����%|	��E�   ��E�   �;|	��E�������E������} v�EP�M�����P�M�Q�]�����j j�M�肹���E�P�M��Q�����R�M��������N����E�M؉H�EP�M�����R��P��|	�;���XZ�M�d�    Y_^[�M�3�������  ;��Z�����]� �   �|	����   �|	_Ptr ���������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��������Iu�E���3�_^[��]������������������������������U����   SVWQ��$����7   ������Y���3ŉE��M�E�P�M������E�P�MQ�UR������R��P�`~	����XZ_^[�M�3��"������   ;��������]� ��   h~	����   t~	_Alval �����������������������������������������������������U����  SVWQ��(����v   ������Y���3ŉE��M�ǅ����    �E�x@ t�E��HE��u��E  �@  �E�   ������P�E��M�B��;��	�����0���������<�����0���Q��<���R�����������t2���  j j�M��׸���E�P��T���Q�M���������������M�������V��h���R�M��~���������P�E��HP�M�I@������H�����h���������T���������H�����(�����(��� t��(���t��(����
  �  �E��@E ��|���P�M��������)����M�+ȉM���|����M����}� vD�E�HPQ�U�Rj������P�M�������������������P�������9E�tǅ(���   �
ǅ(���    ��(�����������������t��������������������������tƅ���� �M��ز���������q�E��HE��uƅ�����M�趲���������O�}� uj j�M�螺���.ƅ�����M�苲���������$ƅ���� �M��t�����������,����M��_���R��P�x�	����XZ_^[�M�3��������  ;��������]Ë�   ��	����   ��	����   ��	_Str _Dest ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�ƅ/��� �E��M�H��/���R�M��E���EP�������_^[���   ;��u�����]� ����������������������������U����   SVWQ��$����7   ������Y���3ŉE��M�M�������M������E�Q�M��j���j�E�Q�M������E��     R��P�t�	����XZ_^[�M�3��������   ;��������]Ð   |�	����   ��	_Alproxy �����������������������������������������������U����   SVWQ��$����7   ������Y���3ŉE��M�M�覫���M��1����E�Q�M�����j�E�Q�M������E��     R��P�T�	����XZ_^[�M�3��+������   ;��������]Ð   \�	����   h�	_Alproxy �����������������������������������������������U����   SVW��@����0   �������EP�MQ����B��0  �у�;��P���_^[���   ;��@�����]��������������������������U����   SVWQ��4����3   ������Y�M��M�{����E_^[���   ;��������]� ����������������������������U����   SVWQ��4����3   ������Y�M��M�	����E_^[���   ;�������]� ����������������������������U���  SVW�������F   ������ǅ8���    �} ��   �E�8 ��   h�  h�a�����Pj�W����������������� t1j �M�����P�������a�����8���P������������������
ǅ����    �E���������8�����t��8���������������   _^[��  ;�������]��������������������������������������������������������������U���  SVW�������F   ������ǅ8���    �} ��   �E�8 ��   h�	  h�a����Pj�7����������������� t1j �M����P�������A�����8���P������襴���������
ǅ����    �E���������8�����t��8�����������~����   _^[��  ;��d�����]��������������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��8 uǅ0���    ��M�����0�����0���_^[��]��������������������������������U����   SVWQ������?   ������Y�M��� ���P�������������P������H������P������E������������P������H������P�E_^[���   ;��%�����]� ��������������������������������������������U����   SVWQ������:   ������Y�M��E���U;Qs�E���Q�E��������
ǅ���    ������U�}� u�E���Q��u�E��9�7������E��E��M;Hs�U��B�M��������
ǅ���    �����_^[���   ;��9�����]� ������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��8 uǅ0���    ��M������0�����0���_^[��]�������������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��0����4   ������Y�M��E��H�9 t�U��B,���0����
ǅ0���    ��0����_^[��]���������������������������U����   SVWQ��0����4   ������Y�M��E��H,����E��H,��E��H�����0����E��H��0������0���_^[��]�������������������������������U����   SVWQ��0����4   ������Y�M��E��H,����E��H,��E��H���0����E��H����E��H���0���_^[��]�����������������������������U����   SVWQ��0����4   ������Y�M��E��H,����E��H,��E��H�����0����E��H��0������0���_^[��]�������������������������������U����   SVWQ��0����4   ������Y�M��M�����;Es�M�聾���E��H;Ms�E��HQ�UR�M������S�E��t;�}s5�E��M;Hs�U��0�����E��H��0�����0���Rj�M�膨����} u
j �M��.����} vǅ0���   �
ǅ0���    ��0���_^[���   ;�������]� �������������������������������������������������������������U����   SVWQ��$����7   ������Y�M��M������E�M��Z����M���+�;E�sǅ$���    ��U���U쉕$�����$����E�E�;Es�E�E�E�_^[���   ;�������]� ������������������������������������U����   SVWQ��4����3   ������Y�M��E����   ��_^[��]������������������������U���   SVWQ�� ����@   ������Y�M��}uǅ ���   �
ǅ ���    �E��� ����HL�E��@E �M��߷���} tJ�   ��tA�E���E�E�E��E���EԋE���EȋE�P�M�Q�U�R�E�P�M�Q�U�R�M������E��M�HP�E����HH�E��@@    _^[��   ;��j�����]� �����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M�H�E��M�H�E��M�H�E��M�H �E��M�H,�E��M�H0_^[��]� ������������������������������U����   SVWQ��4����3   ������Y�M��E����M��A�E����M��A�E����M��A�E����M��A �E���$�M��A,�E���(�M��A0j j �M��ش��j j j �M�����_^[���   ;�������]����������������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ������9   ������Y�M��� ���P�M蟑���M������P�Q�P�Q�@�A_^[���   ;��E�����]� ����������������������������U����   SVWQ��$����7   ������Y�M��E��@0    �E��@    �E��@    �E��@  �E��@   �@    �E��@     �@$    �E��@(    �E��@,    j �M��a���h  h�d�:���Pj��������,�����,��� t��,���������$����
ǅ$���    �E���$����H0_^[���   ;��6�����]����������������������������������������������������������������U����   SVW��@����0   ������E�M�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��M�Җ������t�E��@@    ��E��M�H@�M��Z���_^[���   ;��T�����]� ���������������������������U����   SVWQ��4����3   ������Y�M��} t �M�足��9Er�M�詳���M�A;Ew2����_^[���   ;��������]� �������������������������U����   SVWQ��0����4   ������Y�M��E��M;Hs�U��B;Ewǅ0���   �
ǅ0���    ��0���_^[��]� ����������������������������������U��j�h��d�    PQ��   SVWQ�������@   ������Y���3ŉE�P�E�d�    �e��M�E��U�Q���ǋ�������t  �E��U�Q��螺����t�E��U�Q��舺�����>����E���  �E��U�Q���������  ������P�M��M�J�^���P�������E؍������(����E�    �E��U�Q��������������E���E��U�Q���������x����E������� ����E�P�� ���Q�ܷ�����Ѕ�tj j�E��U�Q��������'�#�E�P���������QjH�M������Ѕ�u���jj�E��U�Q���������	��E�������E������E��U�Q���S�������t��j j�E��U�Q���Y���2�R��P�0�	�����XZ�M�d�    Y_^[�M�3��R�����  ;�������]� ��   8�	����   D�	_Meta ������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��xP t�E��HPQ�������_^[���   ;�������]����������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVW������9   ������M���������uh@c�M胞���� ���P�M����P�M������ ���蹚���EP�M�D����M襚���E_^[���   ;�������]�����������������������������������������U����   SVWQ��0����4   ������Y�M��E��xr�M��QR薴������0�����E�����0�����0���_^[���   ;�������]����������������������������������������U����   SVWQ��0����4   ������Y�M��E��xr�M��QR��������0�����E�����0�����0���_^[���   ;��������]����������������������������������������U����   SVWQ������:   ������Y���3ŉE��M�E�8 tMj�M��Y����E����M���E܋�U܋A��E܃8 t�E܋�    �ދE��A    �M��Y���R��P��	�����XZ_^[�M�3��m������   ;��&�����]ÍI    �	����   (�	_Lock ������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��8 t]�E�����M�E�8 t�E�;M�t�E����M���E�8 uh�   hX`ha臭�����E�M��Q��E��     _^[���   ;��+�����]�����������������������������������������������������U����   SVWQ������:   ������Y���3ŉE��M�j�M�聕���M�讵���E܃}� tN�E܃8 tF�E܋�Q;Ur�E܋�U;Qs�E܋�7����E���E܋�����E܋�����M܋�벍M��]���R��P��	� ���XZ_^[�M�3��q������   ;��*�����]� �   �	����   $�	_Lock ����������������������������������������������������������������������U��j�h��d�    PQ���   SVWQ��$����3   ������Y���3�P�E�d�    �e��M��E�    �E��U�Q���S�������tK�E��U�Q���������t4�E��U�Q��������贕�����uj j�E��U�Q���(�����2�	��E�������E������M�d�    Y_^[���   ;��������]�������������������������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��H �9 t�U��B0���0����
ǅ0���    ��0����_^[��]���������������������������U����   SVWQ��0����4   ������Y�M��E��H0����E��H0��E��H ���0����E��H ����E��H ���0���_^[��]�����������������������������U��j�h �d�    PQ��  SVWQ�������B   ������Y���3�P�E�d�    �e��M�EP������Q�M��������C����E��E�    �E�P�M�QR�E�HQ�M�������-�EP�M�Q������R�M��ە��������j j �g����L�	��E�������E������M������EЋE�x tH�E�HQ�U�BP�M������E�M�@+A��0   ��P�U�BP�����Q�M��`������e���M��w���kE0E܋M�AkE�0E܋M�A�E�M܉H�M�d�    Y_^[��  ;��>�����]� �����������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��n���;Es>�M��������M��\���+�;us�M������M��E���EP�M�����P�M������_^[���   ;��U�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��u����M���D;�u�E��H<Q�U��B8P�M��Q8R�M�褮��_^[���   ;��������]���������������������������U����   SVWQ��4����3   ������Y�M��M�������M���D;�t�M������M��A8�M��l����M��A<�E���EP�M���DQ�U���DR�M�����_^[���   ;��%�����]�����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 tj�E��Q�ΐ�����E��     _^[���   ;�蟼����]�������������������������U����   SVWQ��4����3   ������Y�M��E��8 tj�E��Q�^������E��     _^[���   ;��/�����]�������������������������U����   SVWQ������<   ������Y�M��E��u�y�E��xrp�E��H�M�E���P�����Q�M��-�����������} v �EP�M�Q������P�U���R�������E��H��Q�U�R��#���P�M��������I����E��@   �EP�M��͋��_^[���   ;��G�����]� ��������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x ~�E��HQ�p������$�E��x }�E��H��,�����,���R豟�����E��HQ�;�����_^[���   ;�胺����]���������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x tn�M������E��HQ�U��BP�M��҇���E��M��@+A��0   ��P�U��BP��/���Q�M�賏�����y���E��@    �E��@    �E��@    _^[���   ;�詹����]���������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��xP t�E��HPQ螻����_^[���   ;�������]����������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��E��M��@+A��0   ��_^[��]�������������������U����   SVWQ��4����3   ������Y�M�hm�_���_^[���   ;��������]��������������������������������U����   SVWQ��4����3   ������Y�M�h�m�����_^[���   ;�薷����]��������������������������������U����   SVWQ��4����3   ������Y�M�h m�P���_^[���   ;��6�����]��������������������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q�^�����_^[���   ;��ζ����]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q�������_^[���   ;��n�����]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q螢����_^[���   ;�������]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q�>�����_^[���   ;�讵����]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q�ޡ����_^[���   ;��N�����]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q�~�����_^[���   ;�������]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q������_^[���   ;�莴����]� ���������������������U����   SVWQ��4����3   ������Y�M��EP�M��&x��_^[���   ;��4�����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�M�走��_^[���   ;��Գ����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�M��[���_^[���   ;��t�����]� ���������������������������U����   SVWQ��4����3   ������Y�M�j �EP�J�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M�j �EP�߬����_^[���   ;�貲����]� �������������������������U����   SVWQ��4����3   ������Y�M�j �EP�k�����_^[���   ;��R�����]� �������������������������U����   SVWQ��4����3   ������Y�M��E����M��B��;������_^[���   ;�������]��������������������U����   SVWQ��4����3   ������Y�M��@aPj �MQ�M��v���_^[���   ;�茱����]� �������������������U����   SVWQ��(����6   ������Y�M��M螈��;Es�M��]����M艈��+E�E�E�;Es�E�E�E��@a+H;Mw�M��\����} vT�E��HM�M�j �U�R�M��}������t3�EP�M�X���EP�M��{����M�AP�C������E�P�M��"����E�_^[���   ;�虰����]� ����������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��@a+H;Mw�M��m����} vE�E��HM�M�j �U�R�M��|������t$�EP�MQ�U��BP�M���o���E�P�M��B����E�_^[���   ;�蹯����]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M�h>  h�f�EP�������EP蕜����P�MQ�M�蝶��_^[���   ;��!�����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M��} th*  h�f�EP�������EP�M���n���ȅ�t �EP�M��I����M+�Q�U�R�M��]����n�E��@a+H;Mw�M�辙���} vL�E��HM�M�j �U�R�M���z������t+�EP�MQ�M������U�BP譣�����E�P�M��~���E�_^[���   ;�������]� ��������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��M�ބ��;Es�M�蝤���M�Ʉ��+E�E�E;E�s�E�E�E�;Eu�EE�P�M��?����MQj �M��!����Bj �E�P�M���y���ȅ�t-�E�P�M蜛��EP�M�返��P荢�����E�P�M��l}���E�_^[���   ;�������]� ����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E;@au�M��×��j �EP�M��y���ȅ�t�EP�MQj �M��Xl���EP�M��|���E�_^[���   ;��&�����]� ���������������������������������������������U����   SVWQ��4����3   ������Y�M�h�  h�f�EP�������EP������P�MQ�M��8���_^[���   ;�葫����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��} th  h�f�EP肾�����EP�M��Xk���ȅ�t �EP�M�蹒���M+�Q�U�R�M��S����=j �EP�M��w���ȅ�t%�EP�MQ�M�耒��P�N������EP�M��-{���E�_^[���   ;�褪����]� �����������������������������������������������������������U����   SVW��@����0   ������EP�MQ�UR谖����_^[���   ;�� �����]��������������������������U����   SVW��@����0   ������E�M��_^[��]������������������U����   SVWQ��4����3   ������Y�M��E�P�M��H���P�M�H����E_^[���   ;��x�����]� �������������������������������U����   SVWQ��4����3   ������Y�M��E�P�M��QR�M跾���E_^[���   ;��
�����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E�P�M��QR�M肜���E_^[���   ;�蚨����]� ���������������������������������U����   SVWQ��0����4   ������Y�M��E��8 t�M����0�����E�����0�����0���_^[��]��������������������������������U����   SVWQ��4����3   ������Y�M��M��]���_^[���   ;��ȧ����]������������������U����   SVWQ��0����4   ������Y�M��E��8 uǅ0����a��M��	���H�����0�����0���_^[���   ;��S�����]�����������������������������U����   SVWQ��4����3   ������Y�M��E��M��@+A��0   ��_^[��]�������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��0����4   ������Y�M��E��x8 u�M����0����	�U��0����EP��0���Q�M��Q���_^[���   ;��������]� �����������������������������������U����   SVWQ��4����3   ������Y�M�j �M��v��_^[���   ;�薥����]��������������������������������U����   SVWQ��4����3   ������Y�M��M��C����E��HQ�U��BP�M���r���E��M��Q�P_^[���   ;�������]��������������������������������U����   SVWQ��4����3   ������Y�M�j �EP�M�����_^[���   ;�貤����]� �������������������������U���P  SVWQ�������T   ������Y�M��E���M��A�E��M��P#Qu��   �E��tj j 豜���   �E��M��P#Q��t5j������P�K�����Ph(d������赦��h�O������Q�h����y�E��M��P#Q��t5j������P������PhDd�������o���h�O������Q�"����3j��(���P�е����Ph`d������:���h�O�����Q����_^[��P  ;��l�����]� �����������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��E�E��xP u	�E�    �0�M��h�������u�E�    �E��HPQ�g�������t�E�    jj �M��rr���E�_^[���   ;�艢����]���������������������������������������������������U����   SVWQ��$����7   ������Y�M��EPj0�x�������,�����,��� t�   �u��,���󥋍,�����$����
ǅ$���    _^[���   ;��ۡ����]� ����������������������������������U����   SVW��<����1   ������} u�E��<�����MQ�UR�EP�,p������<�����<���_^[���   ;��T�����]������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M�����_^[���   ;�������]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M��?���_^[���   ;�萠����]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M�����_^[���   ;��0�����]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�ĳ����_^[���   ;��ԟ����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�d�����_^[���   ;��t�����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP������_^[���   ;�������]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP��}������t苈��P�EP�M�g���E������P�EP�M��f���E_^[���   ;�肞����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��E�P�MQ�M�f���E_^[���   ;�������]� ��������������������U����   SVWQ��4����3   ������Y�M��_^[��]���������������������U����   SVWQ��4����3   ������Y�M�2�_^[��]���������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M��E�M��U �E��   ��t	�   �D�B��E����U�
�E ����U �
�E�;Mt�E �;Mt�E��U ��	���3�_^[��]� ������������������������������������������������U����   SVWQ��0����4   ������Y�M��E+E9Es�M��0�����U+U��0�����0���_^[��]� ����������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M��E_^[��]� �����������������U����   SVWQ��4����3   ������Y�M�h
  hb�EP�MQ������h
  hb�EP�"a�����E+EP�MQ�UR��i�����E_^[���   ;�������]� ���������������������������������������������U����   SVWQ��4����3   ������Y�M��E�M��U �E��   ��t	�   �D�B��E����U�
�E ����U �
�E�;Mt�E �;Mt�E��U ��	���3�_^[��]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M��E���P�MQ�c�����_^[���   ;��̙����]� �������������������U����   SVWQ��4����3   ������Y�M�h�	  hb�EP�MQ�F������	�E���E�E;Et�E���P�M�R�Ԉ�����M��ҋE_^[���   ;��3�����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��E���P�MQ�k����_^[���   ;�輘����]� �������������������U����   SVWQ��4����3   ������Y�M�h�	  hb�EP�MQ�6������	�E���E�E;Et�E���P�M�R��j�����M��ҋE_^[���   ;��#�����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��E�M�3�_^[��]� ��������������������������U����   SVWQ��4����3   ������Y�M��E_^[��]� �����������������U����   SVWQ��4����3   ������Y�M�h�	  hb�EP�MQ�������h�	  hb�EP�]�����E+EP�MQ�UR�e�����E_^[���   ;�������]� ���������������������������������������������U����   SVWQ��4����3   ������Y�M��E��H�_^[��]���������������U����   SVWQ��4����3   ������Y�M��E��H�U��B,�	��_^[��]���������������������U����   SVWQ��0����4   ������Y�M��E��x uǅ0���   �
ǅ0���    ��0���_^[��]����������������������������������U����   SVWQ��4����3   ������Y�M��E�P�M��QR�M�����E_^[���   ;��j�����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E�P�M��QR�M�����E_^[���   ;��������]� ���������������������������������U����   SVW��@����0   ��������_^[��]�������������������������U����   SVWQ��4����3   ������Y�M��E��H �U��B0�	��_^[��]���������������������U����   SVW��<����1   ������E�M�;uǅ<���   �
ǅ<���    ��<���_^[��]��������������������U����   SVWQ��0����4   ������Y�M��M�!���P�M���|������t�M��g��;Euǅ0���   �
ǅ0���    ��0���_^[���   ;��o�����]� ��������������������������������������U����   SVWQ��$����7   ������Y�M��EP��MQ��(���R�E���M��B��;��������芉��_^[���   ;�������]� ���������������������������U����   SVWQ��4����3   ������Y�M��E��H;Ms�M�诉���EP�M���b���E�_^[���   ;��n�����]� �������������������������������������U����   SVWQ������9   ������Y�M��E��H;Ms�M��/����E��H+M;Mw�EP�M��ib���F�} v@�M��y��E�E�E��H+M�M��E�+EP�M�MQ�U�R�a�����E�P�M��!b���E�_^[���   ;�蘑����]� �����������������������������������������������U����   SVWQ��0����4   ������Y�M��M��c����tǅ0���   �
ǅ0���    ��0���_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ�� ����8   ������Y���3ŉE��M�E��U�Q���<T����tW�E�P�M��[����M�� �������t4�E��U�Q���T�����c�����uj j�E��U�Q���'����M��]���E�R��P�\�	豣��XZ_^[�M�3��"t�����   ;��ۏ����]�   d�	����   p�	_Ok ������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��H,�+U�E��H,��E��H�U�E��H�_^[��]� ������������������������������U����   SVW��@����0   ��������_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��E��H4Q�M�����E_^[���   ;�莎����]� ���������������������U����   SVWQ��4����3   ������Y�M��E��H0Q�M����E_^[���   ;��.�����]� ���������������������U����   SVWQ��0����4   ������Y�M��M���_����uǅ0���   �
ǅ0���    ��0���_^[���   ;�踍����]����������������������������������U����   SVWQ��4����3   ������Y�M��E��H�_^[��]���������������U����   SVWQ��4����3   ������Y�M��EP�p����P�M��Fg��_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M���M��B��;��N���_^[���   ;��>�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��M��XS���E��M�H8�E��@<    j �M��y���M��A@�E��x8 uj j�M��Ɲ���E��t�E�P�Y����_^[���   ;�茋����]� �����������������������������������U����   SVW��@����0   ��������_^[��]�����������������������U����   SVWQ��0����4   ������Y�M��E�M��Q�B�M#�tǅ0���   �
ǅ0���    ��0���_^[��]� ����������������������������������U����   SVW��<����1   ������E���uǅ<���    ��UR��y������<�����<���_^[���   ;��G�����]���������������������������������U����   SVW��@����0   ��������e��P�EP�M�?W���E_^[���   ;��������]��������������������������U����   SVWQ��4����3   ������Y�M��E�P�g����_^[���   ;�脉����]������������������������������U����   SVWQ��4����3   ������Y�M��E�P�Ջ����_^[���   ;��$�����]������������������������������U����   SVWQ��4����3   ������Y�M����_^[��]��������������������U����   SVWQ��4����3   ������Y�M��UUU_^[��]������������������U����   SVW��@����0   ������M觎��_^[���   ;��M�����]�����������������������U����   SVW��@����0   ������M�r��_^[���   ;��������]�����������������������U����   SVWQ������:   ������Y�M���#���P�M�� �������e���E�}�wǅ���   ��E������������_^[���   ;��s�����]���������������������������������������������U����   SVWQ��(����6   ������Y�M���/���P�M���\����贇��_^[���   ;��������]��������������������U����   SVWQ��$����7   ������Y�M��EP��e�����E�}� t�E쉅$����
ǅ$����c��$���Q�M�>����E_^[���   ;��t�����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��}uh�c�M�č���E���EP�MQ�M��]���E_^[���   ;�������]� ��������������������������U����   SVWQ��$����7   ������Y�M��EP�Y������E�}� t�E쉅$����
ǅ$����c��$���Q�M�����E_^[���   ;��T�����]� �������������������������������������������U����   SVWQ��0����4   ������Y�M��M��aq����0����M��9Y����P�EP��0������0����B��;��Ʉ���E_^[���   ;�趄����]� �����������������������������U����   SVW��<����1   ������} u�E��<�����MQ�UR�EP�]R������<�����<���_^[���   ;��4�����]������������������������������U����   SVWQ��4����3   ������Y�M��xc_^[��]������������������U����   SVWQ��4����3   ������Y�M���c_^[��]������������������U����   SVWQ��4����3   ������Y�M��d_^[��]������������������U����   SVW��8����2   ��������z���M9t�U���<����+�z����uǅ8���   �
ǅ8���    ��8�����<�����<���_^[���   ;��ۂ����]�������������������������������������U����   SVWQ������9   ������Y�M��E��xP u�EP�MQ�UR������E�}� u3��=j�E�P�M��.R���� ���P�M�蓍��P�8e����P�M��b\���� ����D���E�_^[���   ;�������]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M���M��B��;�莁��_^[���   ;��~�����]� �������������������������������������U����  SVWQ������|   ������Y���3ŉE��M�ǅ����    �x��������EP�����Q��n�����Ѕ�t�EP�r�����3  �W�M���g����t8�M���g�����M��G��;�s"�EP��{�����؋M���O����E��  ��E�xP u
�1x����  �M��g���E�x@ uL�E�HPQ�UR�{������P�NB�����ȅ�t�U��������w�������������  �}  �E�   �EP�9{�����E�j j�M��X���E�P��0���Q�M���u�����������M��@W���V��D���R�M���u��������P�E�P�M�Q�U�R�E��HP�M�I@��W����$�����D�����`����0�����`����$������������� ��  �����~������?  �  ��X���P�M��?u�����f����M�+ȉM���X����`���}� vD�E�HPQ�U�Rj��x���P�M��u�����������#���P�j����9E�tǅ���   �
ǅ���    �������o�����������t���������x����`����o�����t�Kv���������M��R����������   �E��@E�E�9E�t�E�������M���Q���������   �}� v�6�M��U���� sj j�M��Y�����u���������M��Q���������w�h�E�HPQ�U�R�@��������t�M�������u�������������������M��VQ���������(�uu���������M��;Q��������������M��&Q��R��P���	�^���XZ_^[�M�3���a�����  ;��}����]� �I    ��	����   ��	����   ��	����   ��	����   ��	_Str _Dest _Src _Ch ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��s��_^[���   ;���{����]� ������������������U����   SVW��$����7   �����󫡀�3ŉE�j j�E�P�M�w���E�E�E�� R��P���	�;���XZ_^[�M�3��_�����   ;��e{����]Ë�   ��	����   ��	f_buf ��������������������������������������������������U����   SVW������9   ������EP�p�����]��EP�p�����]�EP�p�����]�Q�E��$Q�E��$Q�E��$�M�t���E_^[���   ;��z����]��������������������������������������U���  SVW��������   �����󫡀�3ŉE�h�   ��@����MS��jj@j!�M�}G��P��@�����}����@����H��@��������Ѕ�t,j h�e�������V��������P��]������������a����a������jOj ������P�+f����j jP������P��@����u��j j������P��@����tu��������P�������$������̍�����P�S���������?h����������x�����x������l���ǅ`���    ���`�������`�����`���;�l����  ��@���P��L���Q��b������@���P��8���Q�b������@���P��$���Q�b������@���P�����Q�b�������ċ�����������P������H���ԋ�$������(����J��,����B���̋�8������<����A��@����Q���ċ�L������P����P��T����H������i?��P�������!���j j�����P��@�����s�������������P�M�IL���������^;���������RK����@����}���ER��P���	�|���XZ_^[�M�3���[����  ;��w����]ÍI 
   ��	@����   I�	����P   =�	����   1�	����   /�	����,   *�	L���   #�	8���    �	$���   �	���   �	���   �	dummy v3 v2 v1 normal info h n_triangles header_info stl_file ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ������?   ������Y�M��M���<������   �M��5X�����M���<��;�s~�Dm��������EP�����Q�~c�����Ѕ�u;�M��<���   k���P�;z����������EP�����Q�Cc�����Ѕ�t�M��q���EP�\f�����   �   �E��xP t%�l���� ����EP�� ���Q��b�����Ѕ�t	�l���y�w�E��x@ u6�EP��o������/����M��QPR��/���P�F�����ȅ�t�E�:�8�M���;���M���D;�t!�EP�o�����M��AD�M�� >���E���l��_^[���   ;��nt����]� �����������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��zk��_^[���   ;���s����]� ������������������U����   SVWQ��4����3   ������Y�M��E��H0�+U�E��H0��E��H �U�E��H �_^[��]� ������������������������������U����   SVWQ��4����3   ������Y�M��E��H �_^[��]���������������U����   SVWQ��4����3   ������Y�M��E����M��B4��;���r��_^[���   ;��r����]��������������������U����   SVWQ������<   ������Y�M��EP�g����P�M��RJ���ȅ���   �EP�qg�����M�+A��0   ���E�E��M��P;Qu
j�M��M���E��HQ�U��BP�M��#<��kE�0�M�AP�t:����P�U��BP�����Q�M���G������Z���E��H��0�U��J�g�E��M��P;Qu
j�M��M���E��HQ�U��BP�M��;���EP�:����P�M��QR��#���P�M��WG�����Z���E��H��0�U��J_^[���   ;��\q����]� �����������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@8_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U��j�hP�d�    PQ��  SVWQ�������B   ������Y���3ŉE�P�E�d�    �e��M�h�  h�g�EP�6�����E�    �E��@    �@    j�E�P�M��N���M��TN��������   �E�    �EP�MQ�UR�E��U�Q���3�����k���E��U��E�HM��PU��E�H�P�E�;Eu�M�;Mt	�E؃��E��jj�E��U�Q��膁�����	��E�������E�����j �E�P�M��M�J�Z����E䉅�����M���g��������R��P�D�	�؂��XZ�M�d�    Y_^[�M�3��>S����  ;���n����]� ��   L�	����   X�	_Ok ��������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��M��܃����,�����0�����0��� |$	��,��� v�M�����P��r������(�����E����M��B��;���m����(�����(���_^[���   ;���m����]���������������������������������������U����   SVWQ�� ����8   ������Y���3ŉE��M�M��4���M��D;�u!�}u�E�x@ u�E���M�� �E�M�E�xP tS�M���f������tD�EEu�}t�EP�MQ�UR�E�HPQ�d@������u�E�P�M�QPR�@f������t���P���Q�M�<���E�"�M���S���E�P�M�Q�U�BHP�M�p���ER��P���	�V���XZ_^[�M�3���P�����   ;��l����]� �I    ��	����   ��	_Fileposition ��������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M����P���Q�M�;���E_^[���   ;��k����]� �������������������������������U����   SVWQ������<   ������Y���3ŉE��M�M�p���E�U�M�>��+E�U�EԉU؋E�xP tb�M��d������tS�E�P�M�QPR�g`������u<�E�E�tj�E�P�M�Q�U�BPP�F>������u�E�P�M�QPR�"d������t���P���Q�M�:���E�0�M�/���M�AH�M��Q���E�P�M�Q�U�BHP�M�`n���ER��P���	�*~��XZ_^[�M�3��N�����   ;��Tj����]�  �I    ��	����   ��	_Fileposition ��������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M����P���Q�M�g9���E_^[���   ;��i����]�  �������������������������������U����   SVWQ��4����3   ������Y�M��M��A�Q_^[��]��������������U����   SVWQ��(����6   ������Y�M��E�P��/���Q�N����P�M�Z���E_^[���   ;���h����]� ������������������������U����   SVWQ��(����6   ������Y�M��E�P��/���Q�U����P�M��?���E_^[���   ;��ah����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�P�M�@K���E_^[���   ;��h����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�P�M�	O���E_^[���   ;��g����]� ������������������������U����   SVW��@����0   ������EP�M��2���E_^[���   ;��Fg����]��������������������������������U����   SVW��@����0   ������EP�M�'���E_^[���   ;���f����]��������������������������������U����   SVWQ��0����4   ������Y�M��E��xP tF�} u�EEuǅ0���   �
ǅ0���    �MQ��0���R�EP�M��QPR�Bh������t3���j�E��HPQ�M��6���E�_^[���   ;��'f����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ��4����3   ������Y�M��E��H�U��E��H�U��E+E�M��Q,�_^[��]� ��������������������������������U����   SVWQ��4����3   ������Y�M��E��H�U��E��H �U��E+E�M��Q0�_^[��]� ��������������������������������U����   SVWQ��4����3   ������Y�M��} t�EP�M��6��EP�M��X��_^[���   ;��d����]� ������������������������U����   SVWQ��(����6   ������Y�M��M���y����,�����0�����0��� |$	��,��� v�M��?+��P��h������(�����E����M��B��;���c����(�����(���_^[���   ;���c����]���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E���M��B ��;��^c��_^[���   ;��Nc����]� �������������������������������������U����   SVWQ��4����3   ������Y�M�3�3�_^[��]�������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��M��@+A��0   ��_^[��]�������������������U����   SVWQ������=   ������Y�M��M���w����������������� |$	�����v�M���K��P��f����������]�M���/���� ����{Y����,����� ���P��,���Q�O�����Ѕ�t�SY���������M��bq����������������������_^[���   ;��|a����]����������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ������:   ������Y�M��E��xP ti�aX����P�M���M��B��;��`���� ����?X����,����� ���Q��,���R�vN��������u�M��QPR�Nj������}ǅ��������
ǅ���    �����_^[���   ;��>`����]��������������������������������������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVW��@����0   ��������_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��E��@<_^[��]�����������������U����   SVW��@����0   ������E� _^[��]�����������������������U����   SVW��@����0   ������E� _^[��]����������������������U����  SVWQ�� ����x   ������Y���3ŉE��M�M��%����t.�M��%�����M��@��;�s�M��ps��P�4c�����  ��E�xP u
��U���  �M��ZE���E�x@ uM�E� �E�HPQ�U�R�7��������t�M�Q��b������ �����U���� ����� ����L  �G  �M��<n���E�HPQ�D�����E��}��u�eU����(����M��+1����(����	  �E�Pj�M��9���E�P�M�Q�U�R�E�P��@���Q�M��kS�����f�����M���4���V��T���R�M��HS�����of��P�E��HP�M�I@�V����4�����T����>����@����w>����4����� ����� ��� �A  �� ���~�� �����   �&  �E�9E���   ��h���P�M���R������e�����M��4���+u��u���h����>���}� ~$�E����E��M�QPR�E�E��Q�M�����֍E�P�Na������|����M���/����|�����   �1������P�M��?R�����fe���M�+�Qj �M��#M���������=���~�M��}3����s�oj������P�M���Q�����"e��Pj�M�Q�q-�����������?=���E�P�`�����������M��G/���������(�fS���������M��,/���������������M��/��R��P��
�Oo��XZ_^[�M�3���?�����  ;��y[����]Ë�   �
����   
����   
����   
����   	
����   
_Src _Dest _Ch _Str _Ch ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ������:   ������Y�M��E����M��B��;���Y���� ����~Q����,����� ���Q��,���R�G��������t�VQ���������M��n��P�o^��������������_^[���   ;��Y����]��������������������������������������������U����   SVWQ������:   ������Y���3ŉE��M�M��M ����t+�M��A �����M��;��;�s�M��+ ��P��]�����d�b�E���M�B��;���X���E��pP��������M�Q�����R�F��������t�E�����E�P�M��M�B��;��X���E�R��P��
�8l��XZ_^[�M�3��<�����   ;��bX����]ÍI    �
����   �
_Meta ������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��jO��_^[���   ;��W����]���������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M���M��B ��;��ZW��_^[���   ;��JW����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ������9   ������Y�M��� ���P�M��o?��P�;�����E썍 ����9���EP�M���c��_^[���   ;��=V����]� ������������������������������������U����   SVWQ��4����3   ������Y�M����EP�M���M��B ��;���U��_^[���   ;���U����]� ����������������������������U���  SVWQ�������B   ������Y���3ŉE��M�fW�fEȃ} �"  
�} �  �M���j���E؉U܃}� |}�}� vu�E;E�|�M;M�s�E�E؋M�M܋E�P�M��@��P�MQ�J�����E�E�E�E�E؋M�M܉EȉM̋E+E؋MM܉E�M�E�P�M�����   �E���M�B��;��T���E��GL���������M�Q������R�B��������t�E�>�E�P�O�����M��U���U�Eȃ��M̃� �EȉM̋E���M�� �E�M������EȋU�R��P�,
��g��XZ_^[�M�3��W8����  ;��T����]� �I    4
����   @
_Meta ��������������������������������������������������������������������������������������������������������������������������U���  SVWQ�������A   ������Y�M�fW�fE؃} �$  
�} �  �M��@���E�U�}� |}�}� vu�E;E�|�M;M�s�E�E�M�M�E�P�MQ�M���9��P�iH�����E�E�E�E�E�M�M�E؉M܋E+E�MM�E�M�E�P�M��6���   �EP�eW������P�M���M��B��;��}R���� ����J��������� ���Q�����R�H@��������t�4�-�E���E�E؃��M܃� �E؉M܋E���M�� �E�M������E؋U�_^[��  ;��R����]� ����������������������������������������������������������������������������������������������������������U����   SVW��@����0   ��������E�$���E�$��Y����_^[���   ;��CQ����]�����������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��rP����E�P�MQ����B�H�у�;��PP���E�_^[���   ;��=P����]� ������������������������������������U����   SVWQ��4����3   ������Y�M��M���A��_^[���   ;���O����]������������������U����   SVWQ��0����4   ������Y�M��EP�M��`����uǅ0���   �
ǅ0���    ��0���_^[���   ;��dO����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M��y���E��t�E�P��b�����E�_^[���   ;���N����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bx��;��N��_^[���   ;��N����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��PH��;��N��_^[���   ;��N����]� �������������������������������������U����   SVWQ������:   ������Y�M��E��x t�   �E��8 t)��E��Q����B<�H�у�;��M���E��     �E��x tS�E��x t@�E��H��,�����,����� ����� ��� tj�� ����D��������
ǅ���    �E��@    _^[���   ;��M����]���������������������������������������������������������������U����   SVW��@����0   ��������>��_^[���   ;��L����]���������������������U���x  SVW�������^   ������EP���1��P�M���(��j h�r�������t(��j �E�P������Q�M��?%����uǅ����   �
ǅ����    �������������������	4����������t�M�Q���M���3���E�  j�E�P�M��s��j�j��EP�M�Q�M��J��j h�r��������'��j �E�P������Q�M��$����uǅ����   �
ǅ����    �������������������l3����������t�M�Q���M��Q3���E�p  j�E�P�M�����j�j��EP�M�Q�M��J��j h�r�������:'��j �E�P������Q�M��$����uǅ����   �
ǅ����    ��������������������2����������t�M�vP���M��2���E��   j�E�P�M��9��j�j��EP�M�Q�M��nI��j h�r������&��j �E�P�����Q�M��h#����uǅ����   �
ǅ����    ������������������22����������t�M��O���M��2���E�9j�E�P�M����j�j��EP�M�Q�M���H���E�P�M�h&���M���1���ER��P��
�q]��XZ_^[��x  ;��I����]Ë�   �
����   �
����   �
str pos ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���T  SVW�������U   ������EP����-��P�M��%��j h�r�������$��j �E�P������Q�M��o!����uǅ����   �
ǅ����    �������������������90����������t�M��M���M��0���E�p  j�E�P�M����j�j��EP�M�Q�M���F��j h�r�������$��j �E�P������Q�M��� ����uǅ����   �
ǅ����    �������������������/����������t�M�CM���M��/���E��   j�E�P�M����j�j��EP�M�Q�M��;F��j h�r������j#��j �E�P�����Q�M��5 ����uǅ����   �
ǅ����    �������������������.����������t�M�L���M���.���E�9j�E�P�M��l��j�j��EP�M�Q�M��E���E�P�M�5#���M��.���ER��P��
�>Z��XZ_^[��T  ;��rF����]ÍI    �
����   �
����   �
str pos ����������������������������������������������������������������������������������������������������������������������������������������������������������������U���0  SVW�������L   ������EP���*��P�M��"��j h�r�������!��j �E�P������Q�M��_����uǅ����   �
ǅ����    �������������������)-����������t�M��J���M��-���E��   j�E�P�M����j�j��EP�M�Q�M���C��j h�r������� ��j �E�P�����Q�M�������uǅ����   �
ǅ����    ������������������,����������t�M�3J���M��q,���E�9j�E�P�M�����j�j��EP�M�Q�M��.C���E�P�M�� ���M��6,���ER��P�8
��W��XZ_^[��0  ;���C����]�   @
����   \
����   X
str pos ��������������������������������������������������������������������������������������������������������������������������������U���  SVW�������C   ������EP���e(��P�M����j h�r������D��j �E�P�����Q�M������uǅ����   �
ǅ����    �������������������*����������t�M�H���M��*���E�9j�E�P�M��F��j�j��EP�M�Q�M��{A���E�P�M����M��*���ER��P��
�V��XZ_^[��  ;��LB����]Ð   �
����   
����   
str pos ��������������������������������������������������������������������������������������������U����   SVW��@����0   ������EP����&��_^[���   ;��A����]�����������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BT�Ѓ�;���@��_^[���   ;���@����]�������������������������U����   SVW��@����0   �������EP����Q<�B�Ѓ�;��@��_^[���   ;��w@����]���������������������������������U����   SVWQ������9   ������Y�M���EP�MQ�� ���R����P�M����   ��;��@��P�M����� ����(���E_^[���   ;���?����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BH�Ѓ�;��o?��_^[���   ;��_?����]�������������������������U����   SVWQ��$����7   ������Y�M��E��x ufh@r����Ph�j�'������,�����,��� t�MQ��,����}H����$����
ǅ$���    �U���$����B�E��x u3���E��x t&�E��8 tǅ$���   �
ǅ$���    ��$����P��EP����Q<��Ѓ�;��e>���M���E��@   �E��8 tǅ$���   �
ǅ$���    ��$���_^[���   ;��">����]� �������������������������������������������������������������������������U����   SVWQ������?   ������Y�M������P�m)����P�M��b-���������������������_^[���   ;��q=����]���������������������������U����   SVWQ��0����4   ������Y�M��E��@   ����H<��Q��;��=���M���E��8 tǅ0���   �
ǅ0���    ��0���_^[���   ;���<����]���������������������������������U����   SVWQ��4����3   ������Y�M��E��8 u����H��#��EP�M��R����H<�Q�҃�;��Y<��_^[���   ;��I<����]� ��������������������������������U����   SVW��<����1   ������} t�E��<�������������<�����<���Q�UR�EP��3����_^[���   ;��;����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E��x t�   �4�E��x u3��'��E��HQ�U��P����Q<�B�Ѓ�;��,;��_^[���   ;��;����]��������������������������������������U����   SVW������:   ������} u3��   �EP�M������E�    �E�    �E�P�M�Q�M���:����tT�}�t�}�u"�EP�M��V��P�P������t�   �*�$�}�u�EP�M��0#������L����t�   ��3�R��P�&
��M��XZ_^[���   ;��#:����]�   &
����   G&
����   D&
����   @&
dat id browse ����������������������������������������������������������������������������������U���p  SVW�������\   ������ǅ����    j h�r���������P��K�����E��������U!���}� u3���   �E�    �E�P�M��K���E�P�M�Q�M��N9������   �}���   �M��� ���E��}� tF�EP�������>��������Pj������Q�M��y�����������.K����tǅ����   �
ǅ����    ��������������������t�������������� ����������t��������������l ����������t�EԉE�������E�R��P�(
��K��XZ_^[��p  ;��8����]Ë�   $(
����   S(
����   O(
����   H(
browse dat id ��������������������������������������������������������������������������������������������������������������������������U���d  SVW�������Y   ������ǅ����    �} u6j h�r�������[��P��I�����E����������} u3��$  �E�    �EP�M������E�P�M�Q�M��7������   �}���   �M������Eă}� tF�EP�������w<��������Pj������Q�M��C������������H����tǅ����   �
ǅ����    ��������������������t��������������S����������t��������������6����������t�E��E��2�+�}�u%�}� t�EP�M��������dH����t�E��E��������E�R��P��*
�I��XZ_^[��d  ;��5����]ÍI    �*
����   �*
����   �*
����   �*
browse dat id ��������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ���������H<��Q��;��4��_^[���   ;��4����]�������������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;��)4���j�EP�
  ��_^[���   ;��	4����]���������������������������������������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;��i3���j�EP��	  ��_^[���   ;��I3����]���������������������������������������������������U����   SVW��<����1   ������=�� tI�}sǅ<���   �	�E��<�����MQ�UR��<���P����Q���   �Ѓ�;��2���j�EP�	  ��_^[���   ;��2����]�����������������������������������������������U����   SVW��<����1   ������=�� ��   �} tK�}sǅ<���   �	�E��<�����MQ�UR��<���P����Q���   �Ѓ�;���1���[�I�}sǅ<���   �	�E��<�����MQ�UR��<���P����Q���  �Ѓ�;��1����EP�MQ��  ��_^[���   ;��n1����]������������������������������������������������������������������������U����   SVW��4����3   ������} tN�E�E��=$� t"�   k���U�<
�u�E��P�x;�������E�P����Q��Ѓ�;��0��_^[���   ;��0����]�������������������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��80��_^[���   ;��(0����]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;���/��_^[���   ;��/����]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��X/��_^[���   ;��H/����]����������������������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;��.���j�EP�)  ��_^[���   ;��.����]���������������������������������������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;���-���j�EP�i  ��_^[���   ;���-����]���������������������������������������������������U����   SVW��0����4   ������} w�E   �=�� t0��EP�MQ�UR����H���   �҃�;��G-����0����j�EP�  ����0�����0����M��E���th�r����
P�>�����E�_^[���   ;���,����]�����������������������������������������������������������U����   SVW��0����4   ������} w�E   �=�� to�} t0��EP�MQ�UR����H���   �҃�;��Q,����0����.��EP�MQ�UR����H���  �҃�;��!,����0�����0����E��j�EP�  ���E��E���th�r����P�}=�����E�_^[���   ;���+����]������������������������������������������������������������������������U����   SVW��4����3   ������} tN�E�E��=$� t"�   k���U�<
�u�E��P��5�������E�P����Q��Ѓ�;��+��_^[���   ;��+����]�������������������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��*��_^[���   ;��*����]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��(*��_^[���   ;��*����]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��)��_^[���   ;��)����]����������������������������������U����   SVW��4����3   ������}s�E   �E��P�������E��}� u3��:�} t�E��Pj �M�Q������E�� �����E����E��$�   �E�_^[���   ;���(����]��������������������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��(��_^[���   ;��p(����]��������������������������U����   SVW��@����0   �������EP�MQ����B��  �у�;��(��_^[���   ;�� (����]��������������������������U����   SVW��@����0   ���������H��   ��;��'��_^[���   ;��'����]����������������������U����   SVW��@����0   ������} t�   k���U�<
�u�   �3�_^[��]����������������������������U����   SVW��@����0   ������} t!��EP����Q��@  �Ѓ�;���&��_^[���   ;���&����]������������������������U����   SVW��@����0   �������hﾭޡ���H��@  �҃�;��t&��_^[���   ;��d&����]������������������������������U����   SVW��@����0   ������E�8 t��E�Q����B��у�;���%���E�     _^[���   ;���%����]�������������������������������U����   SVW��(����6   ������EP�M��0���EP�M���1���E�P�M����M�����ER��P��:
�!9��XZ_^[���   ;��U%����]Ë�   �:
����   �:
s ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M��Bh��;���$��_^[���   ;��$����]� ����������������������������������U����   SVWQ������9   ������Y�M���EP����Q�M��Bd��;��R$���E�}� u3��s��h�r����P�M��Q����B���   �у�;��$���E��}� u3��4��EP�M��Q�U�R����P�M��Bh��;���#���E�E��  �E�_^[���   ;���#����]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��Bx��;��D#��_^[���   ;��4#����]������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��B��;���"��_^[���   ;��"����]� ����������������������U����   SVW��(����6   �������EP��,���Q����B�H(�у�;��`"��P�M�������,����_
���E_^[���   ;��9"����]�����������������������������������U���  SVW�������`   ������} ��   	�}   @v~j hXs����������Pj0j jj �E�U��4�����n
���^hs���$������P�����P�MQ�"�����������	���������	���E�_  �  �} ��   	�}   v{j h\s�������s���Pj0j jj �E�U�
�3������	���^hs���$������P�����P�MQ��������������������������E��   �~�} |x	�}   vmj h`s�����������Pj0j jj �U�M�X	���^hs���$������P�����P�MQ������������w���������l���E�Lj hds������z���P�EP��,���Q������P�UR�������,����)�����������E_^[�Ā  ;�������]��������������������������������������������������������������������������������������������������������������������������������������������������U���  SVW�������E   �����󫡀�3ŉE��E�E��E�    �E��D�0�Mԃ��MԋE��D�x�Mԃ��M��E�   �	�Eȃ��Eȃ}� |I�E�M������E��E���
}�E���0�MԈD��Uԃ��U���E���7�MԈD��Uԃ��U�먋Eԉ�����������s���"���������D� j �E�P�M�����ER��P��A
�!2��XZ_^[�M�3������  ;��K����]�   �A
����    B
hexstring ��������������������������������������������������������������������������������������U����   SVW��(����6   ��������E P�MQ�UR�EP���E�$��,���Q����B�H$�у�;��v��P�M������,����u���E_^[���   ;��O����]�����������������������������������������U����   SVW��(����6   ������j h�  h(���,���P�M��-������!����,��������(�_^[���   ;�������]�����������������������������U����   SVW��@����0   ������j h�  h(��M�q!���(�_^[���   ;��\����]����������������������U����   SVW��(����6   ������j h�  h(���,���P�M�-�����!����,�������(�_^[���   ;�������]�����������������������������U����   SVW��@����0   ������j h�  h(��M� ���(�_^[���   ;��|����]����������������������U����   SVW��@����0   ������h� �M��0����tj h�  h(��M�.����� ���hHsh(��@�����(�_^[���   ;�������]������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� xs�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E�� xs_^[��]��������������U����   SVWQ��4����3   ������Y�M��M�����E��t�E�P��-�����E�_^[���   ;�������]� ������������������������U����   SVW��@����0   �������EP�MQ����B��x  �у�;����_^[���   ;��p����]��������������������������U����   SVW��@����0   �������EP�MQ����B��p  �у�;����_^[���   ;�� ����]��������������������������U����   SVWQ������=   ������Y�M��E��E�}� tM�E쉅 ����� ������������� t%��j��������������;��y��������
ǅ���    �E�    _^[���   ;��P����]������������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ����B��  �у�;��p��_^[���   ;��`����]��������������������������U����   SVWQ������<   ������Y�M������P����Q�M���   ��;�����P�M� ��������I����E_^[���   ;�������]� ��������������������������������������������U����   SVW��@����0   ���������H��  ��;��l��_^[���   ;��\����]����������������������U����   SVWQ��4����3   ������Y�M�����P��M���$  ��;����_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M�����P��M���(  ��;����_^[���   ;������]������������������������������U����   SVW��@����0   ���������H��d  ��;��,��_^[���   ;������]����������������������U����   SVWQ��4����3   ������Y�M�����P��M���  ��;�����_^[���   ;������]������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��T��_^[���   ;��D����]������������������������������U����   SVW��@����0   �������EP����Q��|  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ����B��t  �у�;��p��_^[���   ;��`����]��������������������������U����   SVWQ��4����3   ������Y�M��M�������E�P����Q$�BD�Ѓ�;�������E�P�MQ����B$�HL�у�;������E�_^[���   ;�������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��5����E�P����Q$�BD�Ѓ�;��J����EP�M�Q����B$�H�у�;��(���E�_^[���   ;������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M������E�P����Q$�BD�Ѓ�;������EP�M�Q����B$�Hd�у�;��x���E�_^[���   ;��e����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M�������E�P����Q$�BD�Ѓ�;������E�_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�BH�Ѓ�;��r���M��}���_^[���   ;��Z����]������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B$�HL�у�;������E�_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B�H�у�;��n���E�_^[���   ;��[����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H<�у�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��0����4   ������Y�M���EP�M�Q����B$�H<�у�;��n����uǅ0���   �
ǅ0���    ��0���_^[���   ;��>����]� �������������������������������������U����   SVW������9   ������EP�M������EP�M�Q����B$�H@�у�;������E�P�M�\���M������ER��P��R
�[!��XZ_^[���   ;������]�   �R
����   �R
fn �������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H@�у�;������E�_^[���   ;�������]� ����������������������������������U����   SVW��@����0   ���������H(��Q��;����_^[���   ;������]�������������������������U����   SVW��@����0   ���������H(����;��0��_^[���   ;�� ����]��������������������������U����   SVW��@����0   �������j j ����H,��҃�;�����_^[���   ;������]�����������������������������������U����   SVW��@����0   ���������H,��Q,��;��_��_^[���   ;��O����]�������������������������U����   SVW��@����0   ���������H���   ��;���
��_^[���   ;���
����]����������������������U����   SVW��@����0   ���������H$��QX��;��
��_^[���   ;��
����]�������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B(�H�у�;��'
��_^[���   ;��
����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H0�у�;��	��_^[���   ;��	����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�B(�Ѓ�;��2	��_^[���   ;��"	����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�Bh�Ѓ�;�����_^[���   ;������]����������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B��;��W��_^[���   ;��G����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P��M��B��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�B�Ѓ�;��r��_^[���   ;��b����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�HL�у�;�����_^[���   ;�������]� �������������������������������������U����   SVW��(����6   �������EP�MQ��,���R����H���  �҃�;��z��P�M������,����y����E_^[���   ;��S����]���������������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��m��_^[���   ;��]����]�����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q$�M��B��;�����_^[���   ;�������]� �����������������������������U����   SVW��@����0   �������E�Q����B(�H�у�;�����E�     _^[���   ;��l����]��������������������������������������U����   SVW��@����0   �������E�Q����B(�H�у�;�����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B,�H�у�;�����E�     _^[���   ;��l����]��������������������������������������U����   SVW��@����0   �������E�Q����B,�H0�у�;�����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;�����E�     _^[���   ;��k����]�������������������������������������U����   SVW��@����0   �������EP����Q$�B\�Ѓ�;����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP����Q�B �Ѓ�;����_^[���   ;������]���������������������������������U����   SVW��@����0   �������EP�MQ����B�H(�у�;��#��_^[���   ;������]�����������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B��  �у�;�� ��_^[���   ;�� ����]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H�Q�҃�;��0 ��_^[���   ;��  ����]��������������������������U����   SVW��@����0   �������EP����Q�B�Ѓ�;������_^[���   ;�������]���������������������������������U���  SVW�������E   ������E�P�M�P���M��������uǅ����    �M������������   j�E�P�_�������u*�E�P�o�������uǅ����    �M��m����������Tj�EP�#�������u*�EP��������uǅ���    �M��1���������ǅ���   �M����������R��P��a
�[��XZ_^[��  ;�������]�   �a
����   �a
parent �����������������������������������������������������������������������������U����   SVW��@����0   �������EP�MQ����B�H�у�;������_^[���   ;��������]�����������������������������U����   SVW��@����0   �������EP����Q��  �Ѓ�;��t���_^[���   ;��d�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��   �Ѓ�;������_^[���   ;��������]����������������������������������U����   SVW��@����0   �������EP�MQ����B�H�у�;�����_^[���   ;��s�����]�����������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;�����_^[���   ;�� �����]��������������������������U����   SVW��@����0   �������EP�MQ����B�H�у�;�����_^[���   ;�������]�����������������������������U����   SVW��@����0   �������EP�MQ�UR����H��  �҃�;��-���_^[���   ;�������]�����������������������U����   SVW������9   �������EP�� ���Q����B���  �у�;�����P�M�U���� ����
����E_^[���   ;�������]��������������������������������U����   SVW��@����0   �������EP����Q��L  �Ѓ�;��4���_^[���   ;��$�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��D  �҃�;�����_^[���   ;�������]�����������������������U���$  SVW�������I   ������ǅ8���    �=�� t!������P����7����8����������������B�����8���������������������������R�M�����8�����t��8����������R�����8�����t��8�����������5����E_^[��$  ;��������]�����������������������������������������������������������U����   SVW������9   ������� ���P����Q���  �Ѓ�;��A���P�M������ ���莿���E_^[���   ;�������]������������������������������������U����   SVW������9   ������� ���P����Q�B$�Ѓ�;�����P�M�L���� ��������E_^[���   ;�������]���������������������������������������U����   SVW��@����0   ������j�EP�g������E_^[���   ;��$�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H�Q�҃�;������_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ�UR����H��H  �҃�;��M���_^[���   ;��=�����]�����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bd��;������_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q$�B`�Ѓ�;��f���_^[���   ;��V�����]� �����������������������������U����   SVWQ������<   ������Y�M���E�P�����Q����B$�H �у�;������P�M����������8����E_^[���   ;��������]� �������������������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��T���_^[���   ;��D�����]������������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B0��;������_^[���   ;��������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��t���_^[���   ;��d�����]������������������������������U����   SVWQ������<   ������Y�M���E�P�����Q����B$�H$�у�;������P�M����������H����E_^[���   ;��������]� �������������������������������������������U����   SVWQ������<   ������Y�M��EP�����Q�M��'������s�������輹���E_^[���   ;��H�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B,�M��P��;������_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��d���_^[���   ;��T�����]������������������������������U����   SVWQ������<   ������Y�M������P����Q,�M��B��;������P�M����������<����E_^[���   ;��������]� �������������������������������U����   SVWQ������<   ������Y�M������P����Q,�M��B<��;��_���P�M����������謷���E_^[���   ;��8�����]� �������������������������������U����   SVWQ��4����3   ������Y�M�����P$��M��Bp��;������_^[���   ;��������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B,��;��g���_^[���   ;��W�����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B��;������_^[���   ;��������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B8��;�����_^[���   ;��w�����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B(��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B��;�����_^[���   ;�������]���������������������������������U����   SVWQ������9   ������Y�M���E�P�� ���Q����B$�H�у�;��+���P�M������ ����*����E_^[���   ;�������]� �������������������������������������������U����   SVWQ������9   ������Y�M���EP�� ���Q����B,�M��P@��;�����P�M������ ��������E_^[���   ;��d�����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H,�Q�҃�;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B4��;��w���_^[���   ;��g�����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B(��;�����_^[���   ;��������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B ��;��'���_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B$��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP����Q(�M����   ��;�����_^[���   ;�������]�( ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR����P(�M��B��;�����_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����;�����_^[���   ;��������]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����   ��;�����_^[���   ;��s�����]� ��������������������������U����   SVWQ��$����7   ������Y�M��E�P�M�良����u3��.�E��tǅ$���   �
ǅ$���    �M��$�����   R��P�ly
����XZ_^[���   ;��������]�    ty
����   �y
c ����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��?���_^[���   ;��/�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P(�M��B��;������_^[���   ;�������]� ����������������������������������U����   SVWQ��0����4   ������Y�M��} t2��EP�M�Q����B �H$�у�;��H�����tǅ0���   �
ǅ0���    ��0���_^[���   ;�������]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�UR����H �QL�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��BX��;��"���_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B`��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��D���_^[���   ;��4�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;������_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;��K���_^[���   ;��;�����]� ����������������������������������U����   SVWQ������?   ������Y�M��M������E�P�M��������uǅ���    �M������������$�E�P�M����ǅ���   �M����������R��P��~
�E���XZ_^[���   ;��y�����]�    �~
����   �~
str ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;������_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��  �у�;��k���_^[���   ;��[�����]� ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B���   �у�;������_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��o���_^[���   ;��_�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bx��;�����_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��0����4   ������Y�M��EP�M��������tE�M��Q�M�������t2�U��0R�M�������t�E��HP�M�������tǅ0���   �
ǅ0���    ��0���_^[���   ;��������]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��O���_^[���   ;��?�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bt��;������_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��o���_^[���   ;��_�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M����   ��;������_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M���  ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��0����4   ������Y�M��EP�M��{�����t2�M��Q�M��h�����t�U��R�M��U�����tǅ0���   �
ǅ0���    ��0���_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��o���_^[���   ;��_�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bh��;�����_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bp��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bx��;��2���_^[���   ;��"�����]� �������������������������U����   SVWQ��0����4   ������Y�M��EP�M��������tE�M��Q�M�������t2�U��R�M��ϧ����t�E��$P�M�輧����tǅ0���   �
ǅ0���    ��0���_^[���   ;��k�����]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;������_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bp��;�����_^[���   ;��r�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B|��;�����_^[���   ;�������]� �������������������������U����   SVWQ��0����4   ������Y�M��EP�M��;�����t2�M��Q�M��(�����t�U��R�M�������tǅ0���   �
ǅ0���    ��0���_^[���   ;��^�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;������_^[���   ;��������]� ����������������������U����   SVWQ������?   ������Y�M��E�    �E�    �E�P�M��&�����u3���   �}� u)������7���P�M����������i����   �   ��h�s����P�M�Q����B���   �у�;������E��}� uj��M�����3��Lj �E�P�M�Q�M�������u�E�P�e�����3��&j �E��P�M�Q�M������E�P�@������   R��P���
�e���XZ_^[���   ;�������]�    ��
����   
����   ��
c len ������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;������_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��_���_^[���   ;��O�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B\��;������_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bd��;�����_^[���   ;��r�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bl��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bt��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bd��;��2���_^[���   ;��"�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bl��;������_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��O���_^[���   ;��?�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;������_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B`��;��r���_^[���   ;��b�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bh��;�����_^[���   ;��������]� �������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;�����_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P(�M��B$��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q�B�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H4�у�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B4��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��/���_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H8�у�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q$�M��Bl��;��B���_^[���   ;��2�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H$�QP�҃�;������_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�HT�у�;��N���_^[���   ;��>�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B��;������_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H�у�;��^���_^[���   ;��N�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H,�у�;������_^[���   ;��������]� �������������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��`���_^[���   ;��P�����]��������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;������_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�����_^[���   ;��o�����]� ����������������������U����   SVWQ��4����3   ������Y�M���j�EP�MQ����B(�M��P��;�����_^[���   ;��������]� �����������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;�����_^[���   ;��}�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;�����_^[���   ;�������]�����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����   ��;�����_^[���   ;�������]� ��������������������������U����   SVWQ��0����4   ������Y�M��} t	ƅ3����ƅ3��� ��3���P�M������_^[���   ;�������]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B,��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B(�M��P ��;��>���_^[���   ;��.�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��} u3��'��EP�M�Q����B �H(�у�;������   _^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��B8��;��1���_^[���   ;��!�����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;������_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��T���_^[���   ;��D�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BT��;��b���_^[���   ;��R�����]� �������������������������U����   SVWQ������<   ������Y�M��� ���P�M����P�M������������ �������������_^[���   ;��ѿ����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BP��;��b���_^[���   ;��R�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��  �у�;�����_^[���   ;��۾����]� ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��   �Ѓ�;��h���_^[���   ;��X�����]����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����   ��;�����_^[���   ;��ӽ����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B(�M��P|��;��n���_^[���   ;��^�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��P\��;�����_^[���   ;��޼����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��������tE�M��Q�M��������t2�U��0R�M��������t�E��HP�M��������tǅ0���   �
ǅ0���    ��0���_^[���   ;�������]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BH��;�袻��_^[���   ;�蒻����]� �������������������������U����   SVWQ��4����3   ������Y�M�����E�$����P(�M��BT��;��*���_^[���   ;�������]� ���������������������������������U����   SVWQ��4����3   ������Y�M�����E�$����P�M��B(��;�誺��_^[���   ;�蚺����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M���  ��;��+���_^[���   ;�������]� ����������������������������������U����   SVWQ��0����4   ������Y�M��E��� �$�M�������tD�M���A�$�M�������t(�U���B�$�M��q�����tǅ0���   �
ǅ0���    ��0���_^[���   ;��Q�����]� ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B<��;��Ҹ��_^[���   ;��¸����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��BH��;��b���_^[���   ;��R�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B@��;�肷��_^[���   ;��r�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��PX��;�����_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$����P�M��B ��;�芶��_^[���   ;��z�����]� ���������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��y�����tE�M��Q�M��f�����t2�U��R�M��S�����t�E��$P�M��@�����tǅ0���   �
ǅ0���    ��0���_^[���   ;�軵����]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BD��;��B���_^[���   ;��2�����]� �������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$����P(�M��BP��;��̴��_^[���   ;�輴����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$����P�M��B$��;��L���_^[���   ;��<�����]� �����������������������������������U����   SVWQ��0����4   ������Y�M��EQ� �$�M��Б����t@�MQ�A�$�M�趑����t&�UQ�B�$�M�蜑����tǅ0���   �
ǅ0���    ��0���_^[���   ;��w�����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B8��;�����_^[���   ;�������]� �������������������������U����   SVWQ������=   ������Y�M�j �M�������E���h�s����P�M�Q����B���   �у�;��q����Eԃ}� uj��M��g���3��dj �E�P�M�Q�M�H����E�P�M�袜����t �M�Q�U�R�M�輹����tǅ���   �
ǅ���    ������E�E�P�z�����E�R��P�d�
����XZ_^[���   ;��ձ����]�    l�
����   x�
mem ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BL��;��"���_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B0��;�貰��_^[���   ;�袰����]� �������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��B<��;��A���_^[���   ;��1�����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;��ѯ��_^[���   ;��������]� ������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��BL��;��b���_^[���   ;��R�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��BD��;�聮��_^[���   ;��q�����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;�����_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B4��;�袭��_^[���   ;�蒭����]� �������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��B@��;��1���_^[���   ;��!�����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;������_^[���   ;�豬����]� ������������������������U���  SVWQ��X����j   ������Y�M��Qq���M���E��8 u��   �EP��l����Ζ��j h�s�������p���P������谖��j j���l���Q������R������P�ח����P������Q襥����P�����R蕥����P�E���
n����tǅX���   �
ǅX���    ��X�����c���������s���������s����������r����������r��������蕓����l�����r����c�����t�E�P�co�����E�_^[�Ĩ  ;��M�����]� ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP趢�����M���E�_^[���   ;�謪����]� �������������������U����   SVWQ��4����3   ������Y�M��E�P�gn����_^[���   ;��T�����]����������������̋�`��`��`��`��`��`��` ��`$��`(��`,��`0��`4��`8��`<��`@��`�������������U����   SVW��@����0   ������EP�M���   Q�UR�+�����_^[���   ;�蛩����]���������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVW��@����0   ������E�M�H4�E�@%d�E�@8�J�E�@<�J�E�@@E�E�@D:^�E�@H�\�E�@L-\�E�@P�s�E�@l@]�E�@X�\�E�@\^�E�@`5^�E�@d]�E�@T"]�E�@h�t�E�@p�]�E�@t]�E�M�H �E�M��E�M�H0�E�M�H(�E�@,    _^[��]����������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U���h  SVW�������Z   ������j h�   ��\���P�+}����j �EP�MQ�UR�EP��\���Q�������E �E�h�   ��\���P�MQ�URj��s����R��P��
�%���XZ_^[��h  ;��Y�����]Ë�   �
\����   ��
np ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M������M���E�_^[���   ;�������]�����������������������������U����   SVWQ��4����3   ������Y�M��E���s� �E���s�@�E�_^[��]���������������������U����   SVWQ��4����3   ������Y�M��E��M��E��@    �E��@    �E�_^[��]� ���������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q������   �H,�у�;��ȡ���E�_^[���   ;�赡����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q������   �H(�у�;��(����E�_^[���   ;�������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��E�@�E�_^[��]� ���������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E��@    �E��@    �E��@    �E�_^[��]�������������������������������U����   SVWQ��4����3   ������Y�M��E�P�������E��     _^[���   ;�蛞����]���������������������U����   SVWQ��4����3   ������Y�M���E�P������   ��Ѓ�;��@���_^[���   ;��0�����]��������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVW��@����0   ������EE_^[��]����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL��  �у�;��K���_^[���   ;��;�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL�QT�҃�;��˜��_^[���   ;�軜����]� ����������������������������������U����   SVW��@����0   �����������   �􋑈   ��;��Y���_^[���   ;��I�����]�����������������������������������U����   SVW��@����0   ���������HL��Q��;�����_^[���   ;��ߛ����]�������������������������U����   SVW��@����0   ���������HL���   ��;�茛��_^[���   ;��|�����]����������������������U����   SVW��@����0   ���������HL����;��0���_^[���   ;�� �����]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL�B\�Ѓ�;�趚��_^[���   ;�覚����]� �����������������������������U����   SVW��@����0   ���������HL��  ��;��L���_^[���   ;��<�����]����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL��   �Ѓ�;��ә��_^[���   ;��Ù����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M��B��;��X���_^[���   ;��H�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�BX�Ѓ�;�����_^[���   ;��Ҙ����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL���   �у�;��k���_^[���   ;��[�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�BP�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ����BL�M���H  ��;��o���_^[���   ;��_�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;�����_^[���   ;��o�����]�������������������������U����   SVW��@����0   �������EP������   ���   �Ѓ�;�����_^[���   ;�������]���������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;�襕���E�     _^[���   ;�茕����]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��%����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;�襔���E�     _^[���   ;�茔����]��������������������������������������U���0  SVWQ�������L   ������Y�M��M��lV��h�  ������诅��P�������y���j �E�P������Q�M���V����uǅ����   �
ǅ����    �������������������[�����������tǅ���    �M��p���������M��st��������M��xp�������R��P���
�@���XZ_^[��0  ;��t�����]Ð   ��
����   ��
dat ��������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B`�Ѓ�;��Ғ��_^[���   ;������]����������������������������U����   SVW��@����0   ���������H�􋑘   ��;��l���_^[���   ;��\�����]����������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B4�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M����   ��;�菑��_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B0�Ѓ�;��"���_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;�諐��_^[���   ;�蛐����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����QL�M���l  ��;��#���_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;�諏��_^[���   ;�蛏����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B,�Ѓ�;��2���_^[���   ;��"�����]����������������������������U����   SVWQ��4����3   ������Y�M���j �E�P����QL�B8�Ѓ�;������_^[���   ;�谎����]��������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M����   ��;��O���_^[���   ;��?�����]� ����������������������U����   SVWQ������:   ������Y�M���EP�M�Q�����R����HL��  �҃�;��Ս��P�M�ċ��������R���E_^[���   ;�讍����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL�Hh�у�;��>���_^[���   ;��.�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL��D  �Ѓ�;�迌��_^[���   ;�诌����]�������������������������U���0  SVWQ�������L   ������Y�M��M��N��h�  ��������}��P���������j �E�P������Q�M��)O����uǅ����   �
ǅ����    ������������������苉����������tǅ���    �M���h���������M��l��������M��h�������R��P���
�p���XZ_^[��0  ;�褋����]Ð   ��
����   ��
dat ��������������������������������������������������������������������U����   SVWQ������:   ������Y�M���EP�M�Q�����R����HL�Q�҃�;������P�M����������*O���E_^[���   ;��ъ����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M���p  ��;��[���_^[���   ;��K�����]� ����������������������������������U���  SVWQ�������F   ������Y�M��M��,L��h�  ������o{��P�������9}��j �E�P������Q�M��L����uǅ����   �
ǅ����    ������������������������������t�M�d���M��Xf���E��M��}z��P�M�����M��:f���ER��P� �
����XZ_^[��  ;��9�����]�    �
����   �
dat ������������������������������������������������������������������������U���  SVWQ�������F   ������Y�M��M���J��h�  ������z��P��������{��j �E�P������Q�M��iK����uǅ����   �
ǅ����    �������������������˅����������t�M�?c���M��e���E��M��-y��P�M趑���M���d���ER��P�P�
赛��XZ_^[��  ;�������]�    X�
����   d�
dat ������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BL�Ѓ�;��?���_^[���   ;��/�����]�������������������������U����   SVW��@����0   ���������H�􋑜   ��;��܆��_^[���   ;��̆����]����������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;��r���_^[���   ;��b�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL��(  �Ѓ�;������_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;�蒅��_^[���   ;�肅����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;��"���_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;�评��_^[���   ;�蟄����]�������������������������U���0  SVWQ�������L   ������Y�M��M��F��h�  ��������u��P�������w��j �E�P������Q�M��G����uǅ����   �
ǅ����    �������������������{�����������tǅ���    �M��`���������M��d��������M��`�������R��P���
�`���XZ_^[��0  ;�蔃����]Ð   ��
����   ��
dat ��������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;�����_^[���   ;��߂����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL�Q@�҃�;��{���_^[���   ;��k�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M����  ��;������_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP������   �M����   ��;�茁��_^[���   ;��|�����]� �����������������������������������U���8  SVWQ�������N   ������Y�M��M��\C��h�  �������r��P�������it��j �E�P������Q�M���C����uǅ����   �
ǅ����    �������������������K~����������t ��s�� ����M��]��݅ �����M���|��ݝ����M��b]��݅���R��P���
�*���XZ_^[��8  ;��^�����]ÍI    ��
����   ��
dat ����������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;����_^[���   ;������]�������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��BP��;��D��_^[���   ;��4����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �B8�Ѓ�;���~��_^[���   ;��~����]�������������������������U���  SVWQ�������F   ������Y�M��M��@��h�  �������o��P�������q��j �E�P������Q�M��9A����uǅ����   �
ǅ����    �������������������{����������t�M�����M���Z���E�,�M��vU���M���P�Q�P�Q�@�A�M��Z���ER��P���
�u���XZ_^[��  ;��}����]�    ��
����   ��
dat ������������������������������������������������������������������������U���  SVWQ�������F   ������Y�M��M��L?��h�  ������n��P�������Yp��j �E�P������Q�M���?����uǅ����   �
ǅ����    �������������������;z����������t�M跁���M��xY���E�,�M��T���M���P�Q�P�Q�@�A�M��JY���ER��P���
����XZ_^[��  ;��I|����]�    ��
����   �
dat ������������������������������������������������������������������������U���  SVWQ�������F   ������Y�M��M���=��h�  ������/m��P��������n��j �E�P������Q�M��y>����uǅ����   �
ǅ����    ��������������������x����������t�M�W����M��X���E�,�M��R���M���P�Q�P�Q�@�A�M���W���ER��P�P�
赎��XZ_^[��  ;���z����]�    X�
����   d�
dat ������������������������������������������������������������������������U���  SVWQ�������F   ������Y�M��M��<��h�  �������k��P�������m��j �E�P������Q�M��=����uǅ����   �
ǅ����    �������������������{w����������t�M��~���M��V���E�,�M��VQ���M���P�Q�P�Q�@�A�M��V���ER��P���
�U���XZ_^[��  ;��y����]�    ��
����   ��
dat ������������������������������������������������������������������������U���0  SVWQ�������L   ������Y�M��M��,;��h�  �������oj��P�������9l��j �E�P������Q�M��;����uǅ����   �
ǅ����    �������������������v����������tǅ���    �M��VU���������M��3Y��������M��8U�������R��P��
� ���XZ_^[��0  ;��4x����]Ð   �
����   �
dat ��������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��B(��;��w��_^[���   ;��w����]������������������������������U����   SVWQ��4����3   ������Y�M�����PL��M���L  ��;��$w��_^[���   ;��w����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �B<�Ѓ�;��v��_^[���   ;��v����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL��  �҃�;��8v��_^[���   ;��(v����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�Bd�Ѓ�;���u��_^[���   ;��u����]����������������������������U���0  SVWQ�������L   ������Y�M��M��7��h�  ��������f��P�������h��j �E�P������Q�M��)8����uǅ����   �
ǅ����    �������������������r����������tǅ���    �M���Q���������M��U��������M��Q�������R��P���
�p���XZ_^[��0  ;��t����]Ð   ��
����   ��
dat ��������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M����   ��;���s��_^[���   ;���s����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL���   �у�;��s��_^[���   ;��{s����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�Bl�Ѓ�;��s��_^[���   ;��s����]����������������������������U���  SVWQ�������F   ������Y�M��M���4��h�  ������/d��P��������e��j �E�P������Q�M��y5����uǅ����   �
ǅ����    ��������������������o����������t�M�Ww���M��O���E�,�M��I���M���P�Q�P�Q�@�A�M���N���ER��P�P�
赅��XZ_^[��  ;���q����]�    X�
����   d�
dat ������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BP�Ѓ�;��?q��_^[���   ;��/q����]�������������������������U����   SVWQ������9   ������Y�M���j �EP�M�Q�� ���R����HL���   �҃�;���p���M���P�Q�P�Q�@�A�E_^[���   ;��p����]� ����������������������������������������������U����   SVWQ������9   ������Y�M���j�EP�M�Q�� ���R����HL���   �҃�;��p���M���P�Q�P�Q�@�A�E_^[���   ;���o����]� ����������������������������������������������U����   SVW��@����0   ������E���M���;��o��_^[���   ;��po����]��������������������������U����   SVW��@����0   �������EP�MQ�U��M�P��;��o��_^[���   ;��o����]���������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�M��M�B��;��n��_^[���   ;��n����]�������������������������U����   SVW��@����0   �������EP�M��M�B��;��;n��_^[���   ;��+n����]���������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����HL���   �҃�;��m��_^[���   ;��m����]� �����������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;��Dm��_^[���   ;��4m����]������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��B<��;���l��_^[���   ;��l����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL�B$�Ѓ�;��Vl��_^[���   ;��Fl����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL��,  �҃�;���k��_^[���   ;���k����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����BL�H(�у�;��Rk��_^[���   ;��Bk����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL�B �Ѓ�;���j��_^[���   ;���j����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL��4  �у�;��[j��_^[���   ;��Kj����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��BH��;���i��_^[���   ;���i����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL���   �҃�;��hi��_^[���   ;��Xi����]� �������������������������������U����   SVWQ��(����6   ������Y�M���E�P����QL���   �Ѓ�;���h���E�}� u)��j �EP�M�Q����BL���   �у�;��h����M��n}��P�M�U��_^[���   ;��h����]� ���������������������������������������������������U���  SVW�������B   ������M��R���M���m���} t�M��Q����u"ǅ����   �M���'���M��?A���������Qj�M��cQ��P�M�}���M��RQ���E�E�E��E�Ph<����-����������M��'���M���@�������R��P���
�[{��XZ_^[��  ;��g����]�   ��
����   ��
����   ��
active mu ������������������������������������������������������������������������������U���  SVW�������B   ������M��NQ���M��l���} t�M��CP����u"ǅ����   �M��&���M���?���������Qj�M��P��P�M�{���M��P���E�E�E��E�Ph=���,����������M��T&���M��?�������R��P���
�z��XZ_^[��  ;��?f����]�    �
����   �
����   �
active mu ������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�����PL��M����  ��;��e��_^[���   ;��te����]������������������������������U����   SVWQ��$����7   ������Y�M��M��C���E�}�t�}�t�}�tǅ$���    �
ǅ$���   ��$���_^[���   ;���d����]���������������������������������U����   SVW��@����0   �������EP�MQ����BL���   �у�;��d��_^[���   ;��pd����]��������������������������U����   SVW��@����0   �������E�Q����B���   �у�;��d���E�     _^[���   ;���c����]�����������������������������������U����   SVW��4����3   �������`^���E��}� u3��a��j �EP�MQ�UR�E�P����Q��h  �Ѓ�;��tc����u+�}� t��E�P����Q@�B�Ѓ�;��Lc���E�    �E�_^[���   ;��2c����]��������������������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;���b��_^[���   ;��b����]������������������������������U����   SVW��@����0   �������j �EPj �MQ�*^����P�UR�EP����Q��h  �Ѓ�;��;b��_^[���   ;��+b����]�������������������������������������U���T  SVWQ�������U   ������Y�M��\���E�}� u3��  �E�    �E�    �E�    �M���#���M��L���E�E��E��E��EPh]  �M��.��j j �E�P�M��J����u��   �M���o���E���E��Eȃ}� ��   �M���D���E��EȉE��E�Ph�   �K'������u�   �}� u�~j �M��~!���Eԃ}� u�i�E�P�M��`P���E�P�Md�����}� t��E�P����Q@�B�Ѓ�;���`���E�    �`����E쉅�����M���9���M���$���������W�}� t��E�P����Q@�B�Ѓ�;��~`���E�    �E�P��c����ǅ����    �M��9���M��$��������R��P� ��s��XZ_^[��T  ;��*`����]� �    ����   3 ����   0 cd ctr �����������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL���   �Ѓ�;��#_��_^[���   ;��_����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����BL��   �у�;��^��_^[���   ;��^����]� ��������������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����Q���   �Ѓ�;��^��_^[���   ;���]����]��������������������������������������U����   SVWQ��4����3   ������Y�M��E��M�H�E��M$�H��hP�
h��
h��
h��
�E��HQ�U R�EP�MQ���E�$�UR�E��HQ�U�R����HL���   �҃�4;��?]��_^[���   ;��/]����]�  ������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR����HL���   �҃�;��\��_^[���   ;��\����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q���   �Ѓ�;��8\��_^[���   ;��(\����]����������������������������������U����   SVWQ��4����3   ������Y�M���j �EP�M�Q����BL�HD�у�;��[��_^[���   ;��[����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�M�Q����BL�HD�у�;��<[��_^[���   ;��,[����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j �EP�M�Q����BL�HH�у�;��Z��_^[���   ;��Z����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�M�Q����BL�HH�у�;��<Z��_^[���   ;��,Z����]� �����������������������������������U���  SVWQ�������B   ������Y�M��EP�������;T��h�  ��$����HK��P������M��j������Q�����R�M��| ��������W���������d6��_^[��  ;��wY����]� ����������������������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;��Y��_^[���   ;���X����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;��X��_^[���   ;��{X����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;��X��_^[���   ;���W����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL�H<�у�;��W��_^[���   ;��~W����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;��W��_^[���   ;���V����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��P0��;��V��_^[���   ;��~V����]� �������������������������������������U���  SVWQ�������B   ������Y�M�j�������oP��h�  ��$����G��P������dI��j������P�����Q�M�����������iS���������2��_^[��  ;���U����]���������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL�Q�҃�;��KU��_^[���   ;��;U����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M���t  ��;���T��_^[���   ;��T����]� ����������������������������������U���  SVWQ�������B   ������Y�M��EP�������M��h�  ��$�����E��P������G��j������Q�����R�M����������Q����������0��_^[��  ;��T����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP��������L��h�  ��$����E��P�������F��j������Q�����R�M��L���������P���������40��_^[��  ;��GS����]� ����������������������������������������������U����   SVW��@����0   �������EP�MQ����BL���   �у�;���R��_^[���   ;���R����]��������������������������U���  SVWQ�������B   ������Y�M��EP��������L��h�  ��$�����C��P������E��j������Q�����R�M����������O���������/��_^[��  ;��R����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����  ��;��Q��_^[���   ;��Q����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����  ��;��Q��_^[���   ;��Q����]� ����������������������������������U���  SVWQ�������B   ������Y�M����E�$�������`R��h�  ��$����B��P�������C��j������P�����Q�M��S���������M���������;-��_^[��  ;��NP����]� �����������������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������H��h�  ��$����XA��P������"C��j������Q�����R�M����������'M���������t,��_^[��  ;��O����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������BG��h�  ��$����@��P������bB��j������Q�����R�M�����������gL���������+��_^[��  ;���N����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������F��h�  ��$�����?��P������A��j������Q�����R�M����������K����������*��_^[��  ;��N����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP��������E��h�  ��$����?��P�������@��j������Q�����R�M��L���������J���������4*��_^[��  ;��GM����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������KG��h�  ��$����X>��P������"@��j������Q�����R�M����������'J���������t)��_^[��  ;��L����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������mF��h�  ��$����=��P������b?��j������Q�����R�M�����������gI���������(��_^[��  ;���K����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL���   �у�;��KK��_^[���   ;��;K����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;���J��_^[���   ;��J����]� ����������������������������������U���  SVWQ�������B   ������Y�M��EP�������B��h�  ��$�����;��P������=��j������Q�����R�M����������G����������&��_^[��  ;��J����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M���P  ��;��I��_^[���   ;��I����]� ����������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�BL�Ѓ�;��"I��_^[���   ;��I����]����������������������������U����   SVW��@����0   ���������HL��@  ��;��H��_^[���   ;��H����]����������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M���T  ��;��OH��_^[���   ;��?H����]� ����������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��j �EP�M�Q������   �H�у�;���G���E�_^[���   ;��G����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��E���P�J����_^[���   ;��AG����]���������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;���F��_^[���   ;���F����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B�Ѓ�;��fF��_^[���   ;��VF����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B�Ѓ�;���E��_^[���   ;���E����]� �����������������������������U����   SVW��@����0   ���������H0�􋑤   ��;��|E��_^[���   ;��lE����]����������������������U����   SVW��@����0   ���������H8����;�� E��_^[���   ;��E����]��������������������������U����   SVW��@����0   ���������H8��Q<��;��D��_^[���   ;��D����]�������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q���  �Ѓ�;��HD��_^[���   ;��8D����]����������������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ����B��  �у� ;��C��_^[���   ;��C����]����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B,�Ѓ�;��6C��_^[���   ;��&C����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B4�Ѓ�;��B��_^[���   ;��B����]� �����������������������������U����   SVW������=   ��������&����u�\h���M��l2���EPh���M���=���EPh���M���=��j �E�PhicMC�����Q��F��������������M��D��R��P�\�U��XZ_^[���   ;���A����]Ë�   d����   pmsg ������������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��l  �҃�;��=A��_^[���   ;��-A����]�����������������������U����   SVW��@����0   �������EP����Q��\  �Ѓ�;���@��_^[���   ;���@����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q0���   �Ѓ�;��_@��_^[���   ;��O@����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B8�HD�у�;���?��_^[���   ;���?����]� �������������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��t?��_^[���   ;��d?����]������������������������������U����   SVW��@����0   �������EP�MQ����B��$  �у�;�� ?��_^[���   ;���>����]��������������������������U����   SVW��@����0   �������EP�MQ����B�Hx�у�;��>��_^[���   ;��>����]�����������������������������U����   SVW��@����0   ���������H���  ��;��,>��_^[���   ;��>����]����������������������U����   SVW��@����0   �������EP���E�$���E�$�MQ����B���   �у�;��=��_^[���   ;��=����]��������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E�P����Q8�B�Ѓ�;��=��_^[���   ;��
=����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H8�Q�҃�;��<��_^[���   ;��<����]� ��������������������������������������U����   SVW��@����0   �������EP����Q��D  �Ѓ�;��<��_^[���   ;��<����]������������������������������U����   SVW��@����0   �������EP����Q��H  �Ѓ�;��;��_^[���   ;��;����]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��-;��_^[���   ;��;����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��:��_^[���   ;��:����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��M:��_^[���   ;��=:����]�����������������������U����   SVW��@����0   ���������H�􋑄   ��;���9��_^[���   ;���9����]����������������������U����   SVW��(����6   �������j �EP�MQ�UR�EP��,���Q����B��t  �у�;��o9��P�M������,����n!���E_^[���   ;��H9����]����������������������������������U����   SVW��@����0   �������E�Q����B0���   �у�;���8���E�     _^[���   ;���8����]�����������������������������������U����   SVW��@����0   �������E�Q����B8�H�у�;��e8���E�     _^[���   ;��L8����]��������������������������������������U����   SVW��@����0   �������E�Q����B8�H@�у�;���7���E�     _^[���   ;���7����]��������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��x  �Ѓ�;��X7��_^[���   ;��H7����]����������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;���6��_^[���   ;���6����]��������������������������U����   SVW��@����0   �������EP�MQ����B�HP�у�;��s6��_^[���   ;��c6����]�����������������������������U����   SVW��@����0   �������EP����Q��,  �Ѓ�;��6��_^[���   ;���5����]������������������������������U����   SVW������<   ������EPj h@t���������P�M�Q�/��������������E�P����Q�B�Ѓ�;��i5���M��t��R��P��*�I��XZ_^[���   ;��@5����]Ð    +����   +s ��������������������������������������������������U����   SVW��4����3   ������j �M�.���E��}� t�E�P��5�����E�P�+����R��P��+�UH��XZ_^[���   ;��4����]Ë�   �+����   �+c ������������������������������������������U����  SVW��(����6  �����󫡀�3ŉE��E�E�E�P�MQh   ������R��<����������PhDt����Q��4  �Ѓ�;���3���E�    R��P��,�tG��XZ_^[�M�3��������  ;��3����]ÍI    �,����   �,t ��������������������������������������������������������������U����   SVW��@����0   �������EP����Q��8  �Ѓ�;��3��_^[���   ;���2����]������������������������������U����   SVW��@����0   ���������H��QH��;��2��_^[���   ;��2����]�������������������������U����   SVW��@����0   ���������H��QD��;��?2��_^[���   ;��/2����]�������������������������U����   SVW��@����0   ���������H��Q<��;���1��_^[���   ;���1����]�������������������������U����   SVW������9   ������EP��MQ�� ���R����H��t  �҃�;��j1�����pB���� ��������E_^[���   ;��E1����]�������������������������������U����   SVW��(����6   �������,���P����Q��  �Ѓ�;���0��P�M�o����,��������E_^[���   ;��0����]������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H�QL�҃�;��P0��_^[���   ;��@0����]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q���  �Ѓ�;���/��_^[���   ;���/����]����������������������������������U����   SVW��(����6   ������M��J5����E�P����Q�B8�Ѓ�;��_/���E�P�M�����M��^���ER��P�1��B��XZ_^[���   ;��'/����]�   1����   $1str ����������������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��.��_^[���   ;��.����]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��-.��_^[���   ;��.����]�����������������������U����   SVW��(����6   �������,���P����Q��  �Ѓ�;���-��P�M�O
����,��������E_^[���   ;��-����]������������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����Q���  �Ѓ�;��-��_^[���   ;��-����]��������������������������������������U����   SVW��@����0   ������E��P��P�M��@Q�U��0R�E�� P�M��Q�UR�EP����Q���   �Ѓ�;��},��_^[���   ;��m,����]���������������������������������������U����   SVW��@����0   ���������H���  ��;��,��_^[���   ;���+����]����������������������U����   SVW��@����0   ���������H�􋑼   ��;��+��_^[���   ;��+����]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B���  �у�;��4+��_^[���   ;��$+����]������������������������������U����   SVW��@����0   �������EP����Q��L  �Ѓ�;���*��_^[���   ;��*����]������������������������������U����   SVW��@����0   ������E�8 t#��E�Q����B��D  �у�;��J*���E�     _^[���   ;��1*����]���������������������������U����   SVW��@����0   �������EP�MQ�UR����H��X  �҃�;���)��_^[���   ;��)����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H��\  �҃�;��])��_^[���   ;��M)����]�����������������������U����   SVW��@����0   �������EP����Q��H  �Ѓ�;���(��_^[���   ;���(����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR����H���  �҃�;��q(��_^[���   ;��a(����]���������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR����H���  �҃�;���'��_^[���   ;���'����]���������������������������U����   SVW��@����0   �������EP�MQ�UR����H��P  �҃�;��}'��_^[���   ;��m'����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H��T  �҃�;��'��_^[���   ;���&����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H��@  �҃�;��&��_^[���   ;��&����]�����������������������U����   SVW��@����0   ���������H���  ��;��<&��_^[���   ;��,&����]����������������������U����   SVW��@����0   ���������H��p  ��;���%��_^[���   ;���%����]����������������������U����   SVW��@����0   �������EP����Q��<  �Ѓ�;��t%��_^[���   ;��d%����]������������������������������U����   SVW��@����0   �������EP�MQ����B�H@�у�;��%��_^[���   ;���$����]�����������������������������U����   SVW��@����0   �������EP�MQ����B��  �у�;��$��_^[���   ;��$����]��������������������������U����   SVW��@����0   �������EP����Q�B�Ѓ�;��'$��_^[���   ;��$����]���������������������������������U����   SVW��@����0   �������EP����Q��\  �Ѓ�;��#��_^[���   ;��#����]������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��D#��_^[���   ;��4#����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQh�2  ����B���   �у�;��"��_^[���   ;��"����]�����������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���   �҃�;��="��_^[���   ;��-"����]�����������������������U����   SVW��@����0   �������EP�MQ����B���   �у�;���!��_^[���   ;���!����]��������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;��d!��_^[���   ;��T!����]������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;��� ��_^[���   ;��� ����]������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;�� ��_^[���   ;��t ����]������������������������������U����   SVW��@����0   �������EP�MQ����B���   �у�;�� ��_^[���   ;��  ����]��������������������������U����   SVW��@����0   �������EP�MQ����B��|  �у�;����_^[���   ;������]��������������������������U����   SVW��@����0   �������EP����Q�B,�Ѓ�;��7��_^[���   ;��'����]���������������������������������U����   SVW��@����0   �������EP����Q��T  �Ѓ�;�����_^[���   ;������]������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��P��_^[���   ;��@����]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��  �Ѓ�;�����_^[���   ;�������]����������������������������������U����   SVW��@����0   ���������H��P  ��;��l��_^[���   ;��\����]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��d  �Ѓ�;�����_^[���   ;�������]����������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVW��@����0   �������EP����Q��,  �Ѓ�;����_^[���   ;�������]������������������������������U����   SVW��@����0   ���������H��<  ��;����_^[���   ;������]����������������������U����   SVW��@����0   ���������H��0  ��;��<��_^[���   ;��,����]����������������������U����   SVW������=   �������f�����u�M� ���E�^h����M���
���EPh����M����j �E�PhicMC�����Q�d�������v��P�M�.���������i����M�������ER��P��E�,.��XZ_^[���   ;��`����]Ð   �E����   �Emsg ����������������������������������������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�����_^[���   ;������]������������������������������U����   SVW������=   �������������u�M�1���E�^h!���M��q	���EPh!���M����j �E�PhicMC�����Q������������P�M���������������M��J����ER��P�XG�,��XZ_^[���   ;�������]Ð   `G����   lGmsg ����������������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��`  �҃�;��=��_^[���   ;��-����]�����������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P����Q���   �Ѓ�;�������u3���E�R��P��H�c+��XZ_^[���   ;������]�   �H����   �H����   �H����   �Hdata sub_id main_id ������������������������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW������9   ������M�������E�P�MQ����B�H|�у�;��k���E�P�M�  ���M������ER��P�J��)��XZ_^[���   ;��3����]�   J����   Jfn �����������������������������������������������������U����   SVW������=   ������j hLGOg���������PhicMC�E�P�^���������������M��b�����u�M������M��W����E��M��A���P�M�\���M��9����ER��P� K�)��XZ_^[���   ;��8����]Ð   K����   Kdat ��������������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P����Q���   �Ѓ�;������u3���E�R��P��K�3(��XZ_^[���   ;��g����]�   �K����   L����   L����   �Kdata sub_id main_id ������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q0���   �Ѓ�;����_^[���   ;������]�������������������������U����   SVW��(����6   �������EP��,���Q����B���  �у�;��=��P�M�������,����<����E_^[���   ;������]��������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B8�H �у�;��>��_^[���   ;��.����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B0���   �у�;����_^[���   ;������]� ��������������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��4��_^[���   ;��$����]������������������������������U����   SVW��$����7   �������EP��(���Q����B���  �у�;����P�M�����(���������E_^[���   ;������]��������������������������������U����   SVW��@����0   ���������H�􋑄  ��;��<��_^[���   ;��,����]����������������������U����   SVW��@����0   �������EP����Q��(  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P����Q���   �Ѓ�;��S����u3���E�R��P�Q��"��XZ_^[���   ;��'����]�   Q����   HQ����   AQ����   <Qdata sub_id main_id ������������������������������������������������U����   SVW��@����0   �������EP�MQ����B��l  �у�;��p��_^[���   ;��`����]��������������������������U����   SVW��(����6   �������EP��,���Q����B���  �у�;�����P�M������,���������E_^[���   ;�������]��������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��t��_^[���   ;��d����]������������������������������U����   SVW��@����0   �������EP�MQ����B��l  �у�;�� ��_^[���   ;�������]��������������������������U����   SVW�� ����8   �������EP��$���Q����B���   �у�;�����U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��U����]�����������������������������������������������U����   SVW��$����7   ������M��;�����E�P����Q���   �Ѓ�;������E�P�M��	���M������ER��P��T�p��XZ_^[���   ;������]Ð   �T����   �Tbc �����������������������������������������������������U����   SVW��@����0   ���������H��`  ��;����_^[���   ;������]����������������������U����   SVW��@����0   �������EP����Q��   �Ѓ�;��
��_^[���   ;��
����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H8�Q$�҃�;��/
��_^[���   ;��
����]� ��������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��	��_^[���   ;��	����]�����������������������U���   SVW�� ����@   �������������u3��^hs���M��j����EPhs���M�����j �E�PhicMC�����Q�����������������������������M��F��������R��P�`W���XZ_^[��   ;�������]Ë�   hW����   tWmsg ��������������������������������������������������������U���   SVW�� ����@   �������������u3��^h#���M��j����EPh#���M�����j �E�PhicMC�����Q�����������������������������M��F��������R��P�`X���XZ_^[��   ;�������]Ë�   hX����   tXmsg ��������������������������������������������������������U����   SVW��@����0   �������EP�MQ����B��h  �у�;��@��_^[���   ;��0����]��������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ����B���  �у� ;��H��_^[���   ;��8����]����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H8�Q(�҃�;�����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H8�Q0�҃�;��K��_^[���   ;��;����]� ����������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���   �҃�;�����_^[���   ;������]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��]��_^[���   ;��M����]�����������������������U����   SVWQ��4����3   ������Y�M���E�P����Q8�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;����_^[���   ;��t����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H8�Q�҃�;����_^[���   ;�������]� ����������������������������������U����   SVW��@����0   �������EP����Q��8  �Ѓ�;����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B8�H8�у�;����_^[���   ;������]� �������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;����_^[���   ;������]�����������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��4��_^[���   ;��$����]������������������������������U����   SVW��(����6   �������EP�MQ�UR��,���P����Q��X  �Ѓ�;�� ��P�M������,����~����E_^[���   ;�� ����]����������������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����Q��h  �Ѓ�;�� ��_^[���   ;��������]��������������������������������������U����   SVW��@����0   ���������H��d  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�MQ����B��@  �у�;��0���_^[���   ;�� �����]��������������������������U����   SVW��@����0   �������EP�MQ����B���   �у�;������_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��P4��;��N���_^[���   ;��>�����]� �������������������������������������U����   SVW��@����0   �������EP����Q�BT�Ѓ�;������_^[���   ;��������]���������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��`���_^[���   ;��P�����]��������������������������U����   SVW��@����0   �������EP����Q��  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��  �҃�;��}���_^[���   ;��m�����]�����������������������U����   SVW��@����0   �������EP����Q�BX�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP����Q�B\�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��4���_^[���   ;��$�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H�Qt�҃�;������_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M����P�U�R����H0���   �҃�(;��'���_^[���   ;�������]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M����P�U�R����H0���   �҃�(;��w���_^[���   ;��g�����]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P����Q0���   �Ѓ�(;������_^[���   ;�������]�$ ����������������������������������U����   SVW��@����0   �������E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR����H���  �҃�$;��5���_^[���   ;��%�����]�������������������������������U����   SVW��@����0   ���������H��Qd��;������_^[���   ;�������]�������������������������U����   SVW��@����0   �������EP����Q�Bl�Ѓ�;��g���_^[���   ;��W�����]���������������������������������U����   SVW��@����0   ���������H��Qh��;������_^[���   ;��������]�������������������������U����   SVW��@����0   �������EP����Q�Bp�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   ���������H��Q`��;��/���_^[���   ;�������]�������������������������U����   SVW��(����6   �������EP�MQ�UR�EP��,���Q����B���  �у�;�����P�M������,����z����E_^[���   ;�������]������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H0���   �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B0���   �у�;�����_^[���   ;�������]� ��������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���   �҃�;�����_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��4����3   ������} 3��^�EP�MQ�UR�EP�t������E��}� |�E��9E�|/�}� }h�s����P������EE�@� �E���E��E�_^[���   ;��������]���������������������������������������U����   SVW��@����0   ������E;Et�&�} t �} t�} t�EP�MQ�UR�!�����_^[���   ;��U�����]�������������������������������U����   SVW��@����0   ������E;Et�&�} t �} t�} t�EP�MQ�UR������_^[���   ;��������]�������������������������������U����   SVWQ��4����3   ������Y�M��M������E�� ht�E�_^[���   ;��l�����]����������������������U����   SVWQ��4����3   ������Y�M��E�� \t�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E���s� �E���s�@�E���s�@�E�_^[��]�������������������������������������U����   SVWQ��4����3   ������Y�M��E�� Lt�E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��E��     �E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E�� Lt��E��HQ����Bl�H�у�;��V���_^[���   ;��F�����]��������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M���j�E��Q����BH��|  �у�;�����_^[���   ;�������]�������������������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P������E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�UR����HH���   �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���   �҃�;��(���_^[���   ;�������]� �������������������������������U����   SVW��@����0   �������EP����QH��Ѓ�;�����_^[���   ;�������]����������������������������������U����   SVW��@����0   �������h�  ����HH��҃�;��H���_^[���   ;��8�����]����������������������������������U����   SVW��4����3   ������h  ��������E��}� u3��tj �EPh�  �M��������u�.�,j �EPh(  �M�������u��j j�M�������E��-�}� t��E�P����Q@�B�Ѓ�;��p����E�    3�_^[���   ;��W�����]�������������������������������������������������U����   SVW��@����0   ���������HH���  ��;������_^[���   ;��������]����������������������U����   SVW��4����3   ������h�  �������E��}� u3��B�EP�MQ�M��κ����u+�}� t��E�P����Q@�B�Ѓ�;��S����E�    �E�_^[���   ;��9�����]���������������������������������������������������U����   SVW��@����0   ���������HH��  ��;������_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�MQ����BH�H�у�;��c���_^[���   ;��S�����]�����������������������������U����   SVW��@����0   �������*E�YE�X�t�,��E�EP�MQ�UR������_^[���   ;��������]����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;��k���_^[���   ;��[�����]� ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����BH��0  �у�;������_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;��k���_^[���   ;��[�����]� ����������������������������������U����   SVW��@����0   �������EP�MQ����BH���  �у�;������_^[���   ;��������]��������������������������U����   SVWQ��4����3   ������Y�M��E�M� +_^[��]� ��������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;��/���_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����HH���  �҃�;�����_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;��/���_^[���   ;�������]�������������������������U����   SVW��@����0   ��������E�$���E�$����s�$�EP�M�0������$�^������$�MQ�M�����_^[���   ;�������]��������������������������������������������U���   SVW�������H   �����󫍍�����ֺ��P�EP�M�Q�M訥�����E�$���E�$���E��$觱�����$���E�$���E�$���E��$�u������$���E�$���E�$���E��$�C������$���������P�EP�M趬��R��P��|����XZ_^[��   ;��J�����]ÍI    �|����   }v ��������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���j �E��Q����BH��|  �у�;�����_^[���   ;�������]�������������������������������������U���D  SVW��������   ������M������E��E�    �M�+����E��E�    �E�    �E�    �E�    �}� u
�   ��  �M�\���=�  �  j h:  �M�����E��M������E�ǅP���    �M������,����M�N����� ����M��������������������E�    �	�E����E��E�;E���   �� ��� ��   j��E�P�� ����J�����t�����t����tek�t��������1���9E�t�k�t��������7���������������;�P���~��������P���k�t������������EԉE��6�E����M�����,�����,����D;Du�Eԃ��E��	�Eԃ��E������}� tj �EP�M�������u
�%  �   �}� tz�M��������tn�M�����;E�ua��hpt� ���%PkM�Q����B���  �у�;��1����E��}� u
��  �  �E�PkM�Q�U�R�M��o���P�Y�������hpt� ���)PkM�Q����B���  �у�;�������E��}� u
�b  �]  �E�PkM�Q�U�R�E�P���������P��� ~K��hpt� ���.P��P�������Q����B���   �у�;��c����E��}� u
��  ��  j��E�P�M蕯����u
��  ��  �}� tj�EP�M��|�����u
�  �  �}� t�M��y����������
ǅ����    �������E��M������E��E�    �E�    �	�E����E��E�;E���  �� ��� ��  j��E�P�� ���蔸����t�����t������  k�t��������w���9E�t�k�t��������8���������ǅ����    ǅ\���    ǅh���    ���h�������h���k�t������������9�h�����  ��h���Pk�t��������I�����u봋�h���Pk�t�������軟����D�����D�������\����U���,��������\�������\�����D�������\����U�����\�������\�����D�������\����U���,����D����\�������\�����D�����   ��\����E�����\�������\�����D�������\����U���,����D����\�������\�����D�����   ��\����E�����\�������\�����D�������\����U���,����D����\�������\�����D�����   ��\����E�����\�������\����=�����\��������������� �v  j�������+���P�E�P������i���ǅ\���    ������;�����|6h�t� ���ZPhpth�h������hpt� ���ZP������������;�����|
�}	  �x	  ��\����M����������}� t3k�����E�kM�M����P�Q�P�Q�P�Q�P�Q�@�Ak�����E�kM�Mȋ��P�Q�P�Q�P�Q�P�Q�@�A��\���;�������   ��\����M���;�������   ��\����M��D���������D�����\����M��T�����8�����8���������������wj�������$�����D�������,����Uԉ�F��D�������,����UԉT�.��D�������,����UԉT���D�������,����UԉT��\�������\��������Eԃ��Eԋ���������������\���;���������������;�����t6h�t� ���wPhpth�h�$�����hpt� ���wP������������;�����t
�  �  ��  �E����M�����,�����,����D;Dtǅ����   �
ǅ����    �������M��}� �  �E�����,���kU�kE�E��
��J�H�J�H�J�H�J�H�R�P�E�����,���kTU��Eԃ�k�M����B�A�B�A�B�A�B�A�R�Q�E�����,���kTU��Eԃ�k�M����B�A�B�A�B�A�B�A�R�Q�}� tB�E�����,���kTU��Eԃ�k�M����B�A�B�A�B�A�B�A�R�Q�E�����,���kU�kE�Eȋ
��J�H�J�H�J�H�J�H�R�P�E�����,����Uԉ�Eԃ��EԋE�����,���kTU�kE�Eȋ
��J�H�J�H�J�H�J�H�R�P�E�����,����UԉT�Eԃ��EԋE�����,���kTU�kE�Eȋ
��J�H�J�H�J�H�J�H�R�P�E�����,����UԉT�Eԃ��Eԃ}� t[�E�����,���kTU�kE�Eȋ
��J�H�J�H�J�H�J�H�R�P�E�����,����UԉT�Eԃ��E�� �E����M�����,�����,����D�D
�0����E�P�s������E�P�g������n  �M�A���=  �[  �M�Ծ���������M覻���������E�    �	�E����E��E�;�����}P�E��������<� u�ۋE��������|� t�E����������EԍP�M���E����������EԍLP��M�뜋�hpt� ��   PkM�Q����B���  �у�;������E��}� u3���  �E�PkM�Q�U�R�E�P�C�������hpt� ��   P��������Q����B���  �у�;����������������� u3��c  ������P��������Q������R������P�������Eԙ+���P�E�P�M�`�����u"�E�P�Ң����������P�â����3��  �M�3����EȋM�6���������ǅ����    ǅ����    �E�    �	�E����E��E�;������)  �E��������<� u��ǅ����    ������������������������M�������;���   ��������;E�}�������������T;U�|hpt� ��   P�������   �����������k�M�k�����Uȋ��A�B�A�B�A�B�A�B�I�J���������������������������Tk�E�k�����Mȋ��P�Q�P�Q�P�Q�P�Q�@�A��������������������E��������|� ��   ��������;E�}�����������;E�|hpt� ��   P�������   �����������k�M�k�����Uȋ��A�B�A�B�A�B�A�B�I�J��������������k�����E�k�����Mȋ��P�Q�P�Q�P�Q�P�Q�@�A���������������E�������������������������E�    �	�E����E��Eԙ+���9E�}#�E��������D�    �E���������   �Ǎ�����P��������E�P�������   �&�E�P�՟�����E�P�ɟ�����E�P轟����3�R��P� ������XZ_^[��D  ;�������]Ë�   (�����   ������   ������   t����   j�����   d�osadr pointsort ngonpointmap opadr sttpadr �W�n�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �������Ef/Ev�E��Ef/Ev�E��E_^[��]�����������������������U����   SVW��@����0   �������EP���E�$�MQ�UR����HH���  �҃�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��5����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��5����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������EP����QH���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��E����E�     _^[���   ;��,�����]��������������������������������������U����   SVW��@����0   �������EP����QH��  �Ѓ�;������_^[���   ;�������]������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��U����E�     _^[���   ;��<�����]��������������������������������������U����   SVW��@����0   �������E P�MQ���E�$�UR�EP�MQ����BH���   �у�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP���E�$�MQ�UR�EP����QH���   �Ѓ�;��+���_^[���   ;�������]�������������������������������������U����   SVW��@����0   �������EP�MQ�UR����HH���  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����BH���  �у�;��4���_^[���   ;��$�����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ������=   ������Y�M��E�    �E�    �E�    �E�8 u*�MQ�M��������uj�M�������uǅ���    �
ǅ���   �U�������E�8 uc�M��Ѽ���} u�EP�MQ�UR�EP�MQ�M�蝜���7�E�E���M��Q����E��}� t�EP�MQ�UR�E�P�MQ�M��f����ыE�8 u�M��<�����tǅ���    �
ǅ���   �M�������E�8 u�M��R����EP�M��-����   �M������} u�EPj �MQ�UR�EP�M������E��uh  �������E�}� u3��^�M����P�M��[����E�E���M��l����E��}� t1�EPj �MQ�U�R�EP�M�胛���Eԃ}� t�E�P�M��&���뾋E�_^[���   ;�������]� �������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��`  �Ѓ�;������_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;��[���_^[���   ;��K�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;��_���_^[���   ;��O�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���E�P����Q@�B,�Ѓ�;��2���_^[���   ;��"�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q@�B,�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��0����4   ������Y�M���j�E�P����QH���   �Ѓ�;��M�����tǅ0���   �
ǅ0���    ��0���_^[���   ;�������]���������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��!��E��HQ����Bl�H�у�;�袿��_^[���   ;�蒿����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;��/���_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR����Hl�Q�҃�;�谾��_^[���   ;�蠾����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;��/���_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��  �҃�;�踽��_^[���   ;�訽����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��  �҃�;��8���_^[���   ;��(�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���j �E�P����QH���   �Ѓ�;�轼��_^[���   ;�譼����]�����������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;��O���_^[���   ;��?�����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��T  �Ѓ�;��߻��_^[���   ;��ϻ����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��  �у�;��k���_^[���   ;��[�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����HH���  �҃�;��ܺ��_^[���   ;��̺����]� �����������������������������������U����   SVWQ��0����4   ������Y�M��E��x ~�   k� �U�
�h�����0����
ǅ0���������0���_^[���   ;��=�����]���������������������������������������U����   SVWQ��(����6   ������Y�M�j h�  �M��&������#����E�M��s������}�u�E���3�_^[���   ;�諹����]�������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��(  �Ѓ�;��?���_^[���   ;��/�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP���E�$�MQ�U�R����HH��0  �҃�;�軸��_^[���   ;�諸����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;��;���_^[���   ;��+�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QH���  �Ѓ�;�賷��_^[���   ;�裷����]� ��������������������������U����   SVWQ������9   ������Y�M��E�P�M�Q�UR�EP�M������E�;Eu�E����E�;Eu�E�����R��P�4������XZ_^[���   ;�������]� �I    <�����   W�����   T�l2 l1 ������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��  �Ѓ�;��_���_^[���   ;��O�����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;�����_^[���   ;��ߵ����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��8  �у�;��{���_^[���   ;��k�����]� ����������������������������������U����   SVWQ������;   ������Y�M���E�P�����Q����BH��\  �у�;�������U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;��K���_^[���   ;��;�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;��ϳ��_^[���   ;�迳����]�������������������������U����   SVWQ��4����3   ������Y�M�h�  �M�����_^[���   ;��c�����]�����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;������_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;�菲��_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR����Hl�Q�҃�;�����_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M�h�  �M��D���_^[���   ;�裱����]�����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��  �Ѓ�;��?���_^[���   ;��/�����]�������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M��Y���_^[���   ;��Ѱ����]���������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��  �Ѓ�;��o���_^[���   ;��_�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���  �҃�;������_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��P  �Ѓ�;�����_^[���   ;��o�����]�������������������������U����   SVWQ��4����3   ������Y�M�����E�$�EP����Q�M����   ��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��4  �Ѓ�;�菮��_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���j�E�P����QH���   �Ѓ�;�����_^[���   ;�������]�����������������������U����   SVWQ��4����3   ������Y�M�h(  �M��T���_^[���   ;�賭����]�����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��,  �҃�;��H���_^[���   ;��8�����]� �������������������������������U����   SVWQ��4����3   ������Y�M�j h(  �M�����_^[���   ;��Ѭ����]���������������������������U���,  SVWQ�������K   ������Y�M��z���E�}� t�} u3���   �M������E��M��k������Eԃ}� u�E���   �E�    �	�Eȃ��EȋM�����9E���   �E�P�M�Q�U�R�E�P�M�1�����u�ȋE��E��	�E����E��E�;E�_�E�����u$�E������M������U��u��D;Du���E���P�M�l���M����T��U��}��t�E�P�M��6q����K����E�R��P�д�8���XZ_^[��,  ;��l�����]� �I    ش����   �����   �b a ������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�    �}u�M��s����E��$�} u�M��#����E���}u�M��Ͼ���E�}� u3���E�P�MQ�M�蝃��_^[���   ;��H�����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��  �у�;��˩��_^[���   ;�軩����]� ����������������������������������U����   SVWQ������;   ������Y�M���EP�MQ���E�$�U�R�����P����QH��  �Ѓ�;��3����M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;��������]� ��������������������������������������������������U����   SVWQ������;   ������Y�M���EP�MQ���E�$�U�R�����P����QH��  �Ѓ�;��c����M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;��+�����]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��\  �Ѓ�;�诧��_^[���   ;�蟧����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���   �҃�;��8���_^[���   ;��(�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;�軦��_^[���   ;�諦����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��p  �҃�;��8���_^[���   ;��(�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��  �҃�;�踥��_^[���   ;�訥����]� �������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��B��;��D���_^[���   ;��4�����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;��Ϥ��_^[���   ;�迤����]�������������������������U����   SVWQ������;   ������Y�M���EP�MQ�����R����P�M����   ��;��U����M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;�������]� ������������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����QH���   �Ѓ�;�蜣��_^[���   ;�茣����]��������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P����QH�B�Ѓ�;�����_^[���   ;�������]� ����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��X  �Ѓ�;�蟢��_^[���   ;�菢����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��,  �Ѓ�;��/���_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M��E���U����q��_^[���   ;��������]� �����������������������U����   SVWQ��4����3   ������Y�M��E�� %�����_^[��]��������������������������U����   SVWQ��0����4   ������Y�M���E��HQ����Bl�H�у�;������} u�   �T��EP�MQ�UR�EP����Ql��Ѓ�;��٠���M��A�E��x tǅ0���   �
ǅ0���    ��0���_^[���   ;�螠����]� �����������������������������������������������������U����   SVWQ��0����4   ������Y�M���EP����QH��x  �Ѓ�;������M���E��8 tǅ0���   �
ǅ0���    ��0���_^[���   ;�������]� ���������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QH��   �Ѓ�;��c���_^[���   ;��S�����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���   �҃�;�����_^[���   ;��؞����]� �������������������������������U����   SVW��@����0   �������E0P�M,Q�U(R�E$P�M Q���E�$���E�$�UR�EP����QH��P  �Ѓ�,;��B���_^[���   ;��2�����]��������������������������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M���������m��_^[���   ;�躝����]��������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;��[���_^[���   ;��K�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E���U���Tz��_^[���   ;��������]� �����������������������U����   SVWQ��0����4   ������Y�M��E����   �uǅ0���   �
ǅ0���    ��0���_^[��]������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H,�у�;�����_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���   �҃�;�舛��_^[���   ;��x�����]� �������������������������������U����   SVW��@����0   ������E;E}�E��E;E~�E��E_^[��]�������������������������������U����   SVWQ��(����6   ������Y�M��EP��x�����E�}� t�EP�M�Q�M��^���E�_^[���   ;�蘚����]� �������������������������������U����   SVWQ��(����6   ������Y�M��EP�MQ��z�����E�}� t�EP�M�Q�M��]���E�_^[���   ;�������]� ���������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;�诙��_^[���   ;�蟙����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��t  �Ѓ�;��?���_^[���   ;��/�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��   �҃�;��Ș��_^[���   ;�踘����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;��K���_^[���   ;��;�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��  �҃�;��ȗ��_^[���   ;�踗����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QH��   �Ѓ�;��C���_^[���   ;��3�����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����BH��|  �у�;�迖��_^[���   ;�诖����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��8  �҃�;��8���_^[���   ;��(�����]� �������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P����QH��t  �Ѓ�;�貕��_^[���   ;�袕����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;��;���_^[���   ;��+�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H@�Q(�҃�;�軔��_^[���   ;�諔����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;��?���_^[���   ;��/�����]�������������������������U����   SVWQ��4����3   ������Y�M���EPj�M�Q����BH���   �у�;��ɓ��_^[���   ;�蹓����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EPj �M�Q����BH���   �у�;��I���_^[���   ;��9�����]� ��������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P����QH��h  �Ѓ�;����_^[���   ;�貒����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;��K���_^[���   ;��;�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��p  �у�;��ˑ��_^[���   ;�軑����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;��K���_^[���   ;��;�����]� ����������������������������������U���   SVWQ�� ����@   ������Y�M�j h�  �M��g���} u�   �uj h�  �M���]���E�}� u3��Y�M���R���EPh�  �M��-]�����E�$h�  �M��Ԡ��j �E�P�M��Q\��ǅ���   �M��T�������R��P����
���XZ_^[��   ;��>�����]� �   �����   �bc �������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��X  �у�;�蛏��_^[���   ;�苏����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��d  �у�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�EP����Q�M��B,��;�蕎��_^[���   ;�腎����]� ����������������������������U����   SVWQ��4����3   ������Y�M���EPj�M�Q����BH���   �у�;�����_^[���   ;��	�����]� ��������������������������������U����   SVWQ������?   ������Y�M��M��[c���E�}� u3��j  �E�    �}u�M��k����E��$�} u�M��z���E���}u�M��ǡ���E��}� u3��  �M��g����E�    �	�Eԃ��EԋM��D���9E���   �E�P�M�M���Eȃ}� u�ϸ   k� �UȋD
P�M��t����t�E���P�M��R���   �� �MȋTR�M�t����t�Eԍ�   Q�M��`R���E����M����U�u�D;Dt.�   ���MȋTR�M�tt����t�Eԍ�   Q�M��R���   k��UȋD
P�M�Et����t�Eԍ�   Q�M���Q��������   _^[���   ;��.�����]� ���������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;��k���_^[���   ;��[�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��PH��;�����_^[���   ;��ފ����]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P����QH��l  �Ѓ�;��b���_^[���   ;��R�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����BH���  �у�;��߉��_^[���   ;��ω����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E�P����QH���  �Ѓ�;��G���_^[���   ;��7�����]� ������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;��ψ��_^[���   ;�迈����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;��_���_^[���   ;��O�����]�������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����QH���  �Ѓ�;�����_^[���   ;��؇����]����������������������������������U����   SVWQ��4����3   ������Y�M���EP���E�$�M�Q����BH���  �у�;��^���_^[���   ;��N�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R����HH���  �҃�0;�贆��_^[���   ;�褆����]�, �������������������������������������������U����   SVW��@����0   �������E0P���E(�$�M$Q�U R�EP�MQ�UR�EP�MQ�UR����HH���  �҃�,;�����_^[���   ;��������]����������������������������������U����   SVWQ��4����3   ������Y�M���E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R����HH���  �҃�0;��d���_^[���   ;��T�����]�, �������������������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����QH���  �Ѓ�;��̄��_^[���   ;�輄����]��������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P����QH��$  �Ѓ�;��B���_^[���   ;��2�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��H  �у�;��˃��_^[���   ;�軃����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��L  �Ѓ�;��O���_^[���   ;��?�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��<  �у�;��ۂ��_^[���   ;��˂����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QH��@  �Ѓ�;��S���_^[���   ;��C�����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;��ہ��_^[���   ;��ˁ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��  �у�;��[���_^[���   ;��K�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��T  �Ѓ�;��߀��_^[���   ;��π����]�������������������������U����   SVWQ��4����3   ������Y�M��qE���M���E�_^[���   ;��s�����]�����������������������������U����   SVWQ��4����3   ������Y�M��E�P�'D�����E��     _^[���   ;�������]���������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]�����������̋�`��`��`��`��`��`��` ��`��������������U����   SVWQ��0����4   ������Y�M��M��������tǅ0���   �
ǅ0���    ��0���_^[���   ;���~����]����������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��M襃���E_^[���   ;���}����]� ����������������������������U����   SVWQ��4����3   ������Y�M��   @_^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U���  SVW��x����b   ������} u3��   j h�   ��<���P�U�����E��\����E��|����E�E��E��<���ǅ@���%d�E�L8�E�*P�E��T�E��M�E��T�E�N�E��8�E��bh�   ��<���P�MQ�URj�iK����R��P�8��̏��XZ_^[�Ĉ  ;�� |����]Ð   @�<����   L�np �����������������������������������������������������������������U����  SVW��(����v   ������ǅ ���    �}( uǅ0���    �M�vc����0����!  �E�    �M轄������  �M��O���M���D������   �EP��H����e���� ���j h�s�������9W���� ���P��l����re���� ���j j���H���Q��l���R������P�f������ ���P������Q�Yt������ ���P������R�Bt������ ��� P�M��\=�����<����uǅ(���   �
ǅ(���    ��(�����?����� ����� t�� ���ߍ������A���� �����t�� ��������A���� �����t�� �����������dA���� �����t�� ������l����GA���� �����t�� ������������a���� �����t�� ������H����A����?�����t(�E(P�M$Q�M��OC��P�UR�EP�MQ�_�����E��M�� ����!�E(P�M$Qj �UR�EP�MQ�_�����E��E�������M�Pa�������R��P�$�����XZ_^[���  ;��y����]ÍI    ,�����   8�icon �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���  SVW��x����b   ������j h�   ��<���P�{P����ǅ\���    �E��|���h�   ��<���P�MQ�URj�&G����R��P�|�艋��XZ_^[�Ĉ  ;��w����]Ë�   ��<����   ��np ���������������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVW��@����0   ������E������� _^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��E��M���j j j �E��Q����B�H�у�;��v���U��B�E�_^[���   ;��yv����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H|�Q�҃�;��v��_^[���   ;���u����]� ����������������������������������U����   SVWQ��(����6   ������Y�M���E�P������   �BX�Ѓ�;��u���E�}� u3���EP�MQ�M��Vs��_^[���   ;��bu����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H|�Q8�҃�;���t��_^[���   ;���t����]� ����������������������������������U����   SVWQ��(����6   ������Y�M���E�P������   �BX�Ѓ�;��ot���E�}� u3���EP�MQ�M��TO��_^[���   ;��Bt����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��9��E��HQ�UR�EP�M��R����H�Q�҃�;��s���M��A�   _^[���   ;��s����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���j j j �E��Q����B�H�у�;��*s���U��B_^[���   ;��s����]������������������������������U����   SVWQ��(����6   ������Y�M�j\�  ���E�}� t	�E�x\ u�<��E�P�M�Q\�҃�;��r���EP�M���b���EP�M��8���EP�M��8���E�_^[���   ;��cr����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�j\��  ���E�}� t	�E�x\ u�0��E�P�M�Q\�҃�;���q���EP�M��)b���EP�M���7���E�_^[���   ;��q����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j\�F  ���E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;��*q���EP�M��ya���E�_^[���   ;��q����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�j\�  ���E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;��p���EP�M��R���E�_^[���   ;��kp����]� ����������������������������������U����   SVWQ������;   ������Y�M�j\�  ���E�}� t	�E�x\ u�0��E�P�M�Q\�҃�;���o���EP������ba��P�M��-`���E�_^[���   ;��o����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j\�V  ���E�}� t	�E�x\ u���E�P�M�Q\�҃�;��:o���E�_^[���   ;��'o����]���������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��(����6   ������Y�M�j`�  ���E�}� t	�E�x` u���E�P�M�Q`�҃�;��jn��_^[���   ;��Zn����]������������������������������������U����   SVWQ��(����6   ������Y�M�jx��  ���E�}� t	�E�xx u�E����E�P�MQ�U�Bx�Ѓ�;���m���E�_^[���   ;���m����]� ���������������������������������������U����   SVWQ������:   ������Y�M�jt�V  ���E�}� t	�E�xt uh���M�`���E�:��EP�M�Q�����R�E�Ht�у�;��m��P�M�`Z��������j���E_^[���   ;���l����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�j|�
  ���E�}� t	�E�x| u3����E�P�MQ�U�B|�Ѓ�;��dl��_^[���   ;��Tl����]� �������������������������������������������U����   SVWQ��0����4   ������Y�M��E�M��;t3���   �E�x uN�E�8 uF�E�x u=�E��x u�M��9 u�U��z uǅ0���   �
ǅ0���    ��0����   �R�E��x uI�E��8 uA�E��x u8�E�x u�M�9 u�U�z uǅ0���   �
ǅ0���    ��0����M�E�x t�E��x t�E�M��P;Qt3��)�E�x t�E��x t�E�M��P;Qt3���   _^[��]� �������������������������������������������������������������������������������������������U����   SVWQ��$����7   ������Y�M�j|�V  ���E�}� t	�E�x| u�   �<��E�P�MQ�U�B|�Ѓ�;��1j����uǅ$���   �
ǅ$���    ��$���_^[���   ;��j����]� ����������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��~����uǅ0���   �
ǅ0���    ��0���_^[���   ;��ti����]� ���������������������������U����   SVWQ��(����6   ������Y�M�jp�  ���E�}� t	�E�xp u������EP�M�Q�U�Bp�Ѓ�;���h��_^[���   ;���h����]� ����������������������������������������U����   SVW��$����7   ������h�   �x  ���E��}� t�E����    u�EP�M�U���E�=��EP�MQ��(���R�E����   �у�;��<h��P�M�}U����(����e���E_^[���   ;��h����]�����������������������������������������������U����   SVWQ������:   ������Y�M�h�   �  ���E�}� t�E샸�    u�E��4��EP�M�Q�����R�E싈�   �у�;��sg���������d���E�_^[���   ;��Ug����]� ��������������������������������������������U����   SVW��4����3   ������j��  ���E��}� t	�E��x u3���E���H��;���f��_^[���   ;���f����]������������������������������U����   SVWQ������?   ������Y�M�h�   �c  ���E�}� t�E샸�    uj �������W��P�M�Y���E�9��EP�����Q�U�M����   ��;��!f��P�M�bS��������c���E_^[���   ;���e����]� �������������������������������������������������U����   SVWQ��(����6   ������Y�M�j<�  ���E�}� t	�E�x< u���EP�M�Q�U�B<�Ѓ�;��fe��_^[���   ;��Ve����]� �����������������������������U����   SVWQ��(����6   ������Y�M�h�   ��  ���E�}� t�E샸�    u���EP�U�M����   ��;���d��_^[���   ;���d����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S  ���E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��'d��_^[���   ;��d����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�j4�  ���E�}� t	�E�x4 u3����E�P�M�Q4�҃�;��c��_^[���   ;��xc����]����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �  ���E�}� t�E샸�    u3����E�M����   ��;���b��_^[���   ;���b����]���������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s   ���E�}� u3��'��EP�MQ�UR�E�P�M싑�   �҃�;��Ob��_^[���   ;��?b����]� ��������������������������������������U����   SVW��@����0   ������h���EPhD �G����_^[���   ;���a����]�������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u3����EP�U�M����   ��;��Oa��_^[���   ;��?a����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�jD��������E�}� t	�E�xD u3����E�P�M�QD�҃�;��`��_^[���   ;��`����]����������������������������������U����   SVWQ��(����6   ������Y�M�jL�F������E�}� u3����EP�M�Q�U�BL�Ѓ�;��-`��_^[���   ;��`����]� ������������������������������������U����   SVW������9   ������h�   �������E��}� u�M�e���E�9��EP�� ���Q�U����   �Ѓ�;��_��P�M�<���� ����G���E_^[���   ;��i_����]���������������������������������������������������U����   SVW��4����3   ������j��������E��}� t	�E��x u3�� ��EP�MQ�UR�E��H�у�;���^��_^[���   ;���^����]�������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��7^��_^[���   ;��'^����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�U�M����   ��;��]��_^[���   ;��]����]� ��������������������������������������U����   SVW��4����3   ������E�8 u�?j�������E��}� t	�E��x u�!��EP�M��Q�҃�;���\���E�     _^[���   ;���\����]��������������������������������������U����   SVWQ��(����6   ������Y�M�jH�v������E�}� u���EP�M�Q�U�BH�Ѓ�;��_\��_^[���   ;��O\����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M��E�    �	�E���E�E�P�M��"0���8 t��E�_^[���   ;���[����]����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� u�'��EP�MQ�UR�E�P�M싑�   �҃�;��A[��_^[���   ;��1[����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�j$��������E�}� t	�E�x$ u3����E�P�M�Q$�҃�;��Z��_^[���   ;��Z����]����������������������������������U����   SVWQ������9   ������Y�M�h�   �3������E�}� t�E샸�    u3����E�M����   ��;��Z���E��E�_^[���   ;���Y����]���������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� u3����EP�M�Q�U싂�   �Ѓ�;��wY��_^[���   ;��gY����]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� u3����EP�M�Q�U싂�   �Ѓ�;���X��_^[���   ;���X����]� ������������������������������U����   SVWQ��(����6   ������Y�M�j8�v������E�}� t	�E�x8 u3��(��EP�MQ�UR�EP�M�Q�U�B8�Ѓ�;��HX��_^[���   ;��8X����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� u3����EP�M�Q�U싂�   �Ѓ�;��W��_^[���   ;��W����]� ������������������������������U����   SVWQ��(����6   ������Y�M�j(�6������E�}� t	�E�x( u3��$��EP�MQ�UR�E�P�M�Q(�҃�;��W��_^[���   ;���V����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j,�������E�}� t	�E�x, u3�� ��EP�MQ�U�R�E�H,�у�;��pV��_^[���   ;��`V����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�jP��������E�}� u3�� ��EP�MQ�U�R�E�HP�у�;���U��_^[���   ;���U����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�jT�f������E�}� u3����E�P�M�QT�҃�;��QU��_^[���   ;��AU����]���������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� u3��/��EP�MQ�UR�EP�MQ�U�R�E싈�   �у�;��T��_^[���   ;��T����]� ����������������������������������������������U����   SVWQ��$����7   ������Y�M��E�    �	�E���E�E�P�M��r(���8 t(�E�P�M�a(��P�M�Q�M��T(������`����t�뾃} t�E�M��}� ~�E�P�M��%(���8 uǅ$���   �
ǅ$���    ��$���_^[���   ;��S����]� �����������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j�6������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;��S��_^[���   ;��S����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;��tR��_^[���   ;��dR����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M��} u3��@j��������E�}� t	�E�x u3�� ��EP�MQ�U�R�E�H�у�;���Q��_^[���   ;��Q����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�jl�F������E�}� t	�E�xl u���E�P�M�Ql�҃�;��*Q��_^[���   ;��Q����]������������������������������������U����   SVWQ��(����6   ������Y�M�jh�������E�}� t	�E�xh u���EP�M�Q�U�Bh�Ѓ�;��P��_^[���   ;��P����]� �����������������������������U����   SVWQ��(����6   ������Y�M�h�   �#������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;���O��_^[���   ;���O����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�U�M����   ��;��_O��_^[���   ;��OO����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��N��_^[���   ;��N����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�jd�6������E�}� t	�E�xd u���EP�M�Q�U�Bd�Ѓ�;��N��_^[���   ;��N����]� �����������������������������U����   SVWQ��(����6   ������Y�M�j(�������E�}� t	�E�x0 u3��$��EP�MQ�UR�E�P�M�Q0�҃�;��|M��_^[���   ;��lM����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�jX�������E�}� u���EP�M�Q�U�BX�Ѓ�;���L��_^[���   ;���L����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j �v������E�}� t	�E�x  u3����E�P�M�Q �҃�;��XL��_^[���   ;��HL����]����������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��K��_^[���   ;��K����]� ����������������������������������U����   SVW��<����1   ������E��<�����<���t��E����E����   _^[��]� ��������������������������������U����   SVW������:   ������E�����������������������q  ������$���   �]  ���������=����   �EP�K����=�2  }
������&  �} u
������  h�t�$���Ph�j�%������ ����� ��� t�� ����G%��������
ǅ���    ���������=�� t�EP����
'���   �   �EP�MQ�P������u����   �   �|��I���u��������u\�6���	���=�� t?�����8�����8�����,�����,��� tj��,����E@��������
ǅ���    ���    �   ����_^[���   ;��LI����]Ðz[bp�8����������������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��M��#���E�    �	�E���E�}�}�E�M��D�    ��E�_^[���   ;��MH����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �M��A    �U��B    �E��@    �E��@    �E�_^[��]�����������������������������������������U����   SVWQ��4����3   ������Y�M��M����A���M��:L���E�_^[���   ;��JG����]��������������������U����   SVWQ��4����3   ������Y�M��M��i��_^[���   ;���F����]������������������U����   SVWQ��4����3   ������Y�M��M��I���M�������_^[���   ;��F����]�����������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B��(  �у�;��;F���E�_^[���   ;��(F����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B��,  �у�;��E��_^[���   ;��E����]� ����������������������������������U����   SVWQ��0����4   ������Y�M���E�P�MQ����B��,  �у�;��;E����uǅ0���   �
ǅ0���    ��0���_^[���   ;��E����]� ����������������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVWQ��4����3   ������Y�M��M��Y���E��t�E�P�DX�����E�_^[���   ;��QD����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H�Q@�҃�;���C��_^[���   ;���C����]� ����������������������������������U����   SVW��@����0   ���������H����;��C��_^[���   ;��pC����]��������������������������U����   SVW��@����0   ���������H���   ��;��C��_^[���   ;��C����]����������������������U����   SVW��@����0   ���������H��   ��;��B��_^[���   ;��B����]����������������������U����   SVW��@����0   ���������H��\  ��;��\B��_^[���   ;��LB����]����������������������U����   SVW��0����4   ������hHu�(���Ph�h�   �"������8�����8��� t��8����LN����0����
ǅ0���    ��0���_^[���   ;��A����]���������������������������������������������U����   SVW��@����0   ���������H����;��PA��_^[���   ;��@A����]��������������������������U����   SVWQ��4����3   ������Y�M��EP�M���U��_^[���   ;���@����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�M��U��_^[���   ;��@����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M�����xX u�'��EP�M��~�����M��t���H �WX��;��	@��_^[���   ;���?����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��������M������H �WH��;��?��_^[���   ;��y?����]� ��������������������������������U����   SVWQ��4����3   ������Y�M��M�����xT u����+��EP�MQ�M��g�����M��]���H �WT��;���>��_^[���   ;���>����]� �����������������������������������������U���  SVWQ�������C   ������Y�M��} t<�M��� ����E�P�M��� �����M��� ���H �WL��;��[>���M��M�����} t?�������
D��P�M��)���������<&���M��} ���@@�EЃ}� t�E�P�M�)��R��P�T"�Q��XZ_^[��  ;���=����]� �I    \"����   h"bc ���������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M������xL u3��/��EP�MQ�UR�M��������M������H �GL��;��=��_^[���   ;��=����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��M������x` u� }  �'��EP�M���������M�������H �W`��;��<��_^[���   ;��t<����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��M��t����xH u3��#�M��b������M��X������H �FH��;���;��_^[���   ;���;����]�������������������������������������U����   SVWQ��4����3   ������Y�M��M�������xX u����'��EP�M���������M�������H �WX��;��V;��_^[���   ;��F;����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��F������M��<����H �G@��;���:��_^[���   ;���:����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��������M������H �GD��;��A:��_^[���   ;��1:����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��M��4����xP u����3��EP�MQ�UR�EP�M��������M������H �WP��;��9��_^[���   ;��9����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��M������xP u������;��EP�MQ�UR�EP�MQ�UR�M��e������M��[����H �GP��;���8��_^[���   ;���8����]� ���������������������������������������U����   SVWQ��$����7   ������Y�M�j�EP��B������tǅ$���   �
ǅ$���    ��$���Q�M���"���E�M���;E��M�"C��;E�~������3��EP�MQ�UR�EP�M��w������M��m����H �WD��;��8��_^[���   ;���7����]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�������xT u������+��EP�MQ�M���������M������H �WT��;��P7��_^[���   ;��@7����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��l  �у�;���6��_^[���   ;��6����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H�Q�҃�;��K6��_^[���   ;��;6����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��@����P�M������Pj j �E�P����Q�B4�Ѓ� ;��5��_^[���   ;��5����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q����B�H4�у� ;��5��_^[���   ;��5����]� �����������������������������U����   SVWQ��4����3   ������Y�M��M��I���M��9��_^[���   ;��4����]��������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��B4��_^[���   ;��24����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H��h  �҃�;��3��_^[���   ;��3����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H���   �҃�;��,3��_^[���   ;��3����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�H\�у�;��2��_^[���   ;��2����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��} t�M�����0����
ǅ0���    ��0���P�M�Q����B��8  �у�;��2��_^[���   ;���1����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B �Ѓ�;��1��_^[���   ;��r1����]����������������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��1����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;���0����]������������������U����   SVW��@����0   �������E�Q����B�H�у�;��u0���E�     _^[���   ;��\0����]��������������������������������������U����   SVW��@����0   �������E�Q����B���   �у�;���/���E�     _^[���   ;���/����]�����������������������������������U����   SVW��@����0   �������E�Q����B��$  �у�;��r/���E�     _^[���   ;��Y/����]�����������������������������������U����   SVW��@����0   �������E�Q����B��`  �у�;���.���E�     _^[���   ;���.����]�����������������������������������U����   SVW��$����7   ������E�8 t?�E���8�����8�����,�����,��� tj��,����s����$����
ǅ$���    �E�     _^[���   ;��5.����]�����������������������������������������������U����   SVW��@����0   �������E�Q����B�H�у�;���-���E�     _^[���   ;��-����]��������������������������������������U����   SVW��@����0   �������E�Q����B�H�у�;��E-���E�     _^[���   ;��,-����]��������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t j j j�E���P�M��	����E��     �E��x` t�E���`P������_^[���   ;��,����]������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q���   �Ѓ�;��,��_^[���   ;��,����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��+��_^[���   ;��+����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��B+��_^[���   ;��2+����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�BP�Ѓ�;���*��_^[���   ;���*����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�HT�у�;��^*��_^[���   ;��N*����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�HT�у�;���)��_^[���   ;���)����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��b)��_^[���   ;��R)����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B�HX�у�;���(��_^[���   ;���(����]� �������������������������U����   SVWQ������<   ������Y�M���h�  �E�P�� ���Q����B���   �у�;��c(�����&	��������� ����(�������_^[���   ;��5(����]�����������������������������������������������U����   SVWQ������9   ������Y�M���EP�MQ�U�R�� ���P����Q���   �Ѓ�;��'��P�M������ ����y���E_^[���   ;��'����]� ��������������������������������U����   SVW��@����0   ���������H��t  ��;��,'��_^[���   ;��'����]����������������������U����   SVW��@����0   ���������H��4  ��;���&��_^[���   ;��&����]����������������������U����   SVW��@����0   ���������H��p  ��;��l&��_^[���   ;��\&����]����������������������U����   SVW��@����0   ���������H��0  ��;��&��_^[���   ;���%����]����������������������U����   SVWQ������9   ������Y�M���EP�M�Q�� ���R����H��L  �҃�;��%��P�M�#���� �������E_^[���   ;��n%����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��} t�E�M��Ap� �E��xd t�E��@h��E��x|u�   �3�_^[��]� ����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�BL�Ѓ�;��$��_^[���   ;��r$����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�BL�Ѓ�;��$��_^[���   ;��$����]����������������������������U����   SVWQ������<   ������Y�M��M�+3���M��r�����uhHu�0���P�25����3��   �E�    ��E�P�M�Q�UR�E�P����Q���   �Ѓ�;��[#����u3��M�E�    �	�Eԃ��EԋE�;E�}"�EԋM��<� u��EԋM���R�M�����͍E�P�������   R��P�T=�6��XZ_^[���   ;���"����]�    \=����   x=����   t=arr count ����������������������������������������������������������������������������������U����   SVWQ������<   ������Y�M��M������M��������uhHu�4���P�3����3��   �E�    ��E�P�M�Q�UR�E�P����Q���   �Ѓ�;���!����u3��i�}� u3��_�E�    �	�Eԃ��EԋE�;E�}4�EԋM��<� t�EԋM����W�����u�ϋEԋM���R�M����뻍E�P��������   R��P��>�5��XZ_^[���   ;��I!����]�    �>����   ?����   ?arr count ��������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�����P��M���|  ��;�� ��_^[���   ;��t ����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q��T  �Ѓ�;�� ��_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q�B�Ѓ�;����_^[���   ;������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B���   �у�;����_^[���   ;�������]� ��������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B��   �у�;����_^[���   ;��t����]������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@`    �E��@d    �E��@h    �E���s�@p�E��@x�����E��@|   _^[��]��������������������������������������������U����   SVW�� ����8   ������M�����E�P�MQ�A*������t�}� u3���E�P�M�Q�U�R�E�P�M�����R��P�C�1��XZ_^[���   ;��6����]ÍI    C����   Cdat ����������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q��P  �Ѓ�;����_^[���   ;������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�Bh�Ѓ�;��2��_^[���   ;��"����]����������������������������U����   SVWQ��4����3   ������Y�M��E��8 thHu�,���P�^-�����E��x` thHu�,���P�?-�����M��,����M��p ���E�P�M���dQ�U��BxP�MQ�U���`R�������M��A|�E��x|u�E��8 u>�E��8 u�E��x|u
�E��@|�����E��     �E���`P�'������E��@|�   �E��xd ��   �E���pP�M���hQ�UR�.������u0�E��@h    �E���s�@phHu�,���P�Z,�����EP�M�������j j j�E���P�M��	������U��B|�E��x|t�M������E��@|��E��@x�����E��@|_^[���   ;��Y����]� ����������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q����B�H�у� ;����_^[���   ;��v����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��<  �у�;����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q��@  �Ѓ�;����_^[���   ;��s����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H��d  �҃�;�����_^[���   ;�������]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E��xd u�E��@`�}�E��M;Hxu�E��@`�j�EP�M��Q`Rj�E���P�M��	�����U��B|�E��x|u �E��M�Hx�} t	�E�    �E��@`��E��@x�����} t�E�M��Q|�3�_^[���   ;������]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�HD�у�;��~��_^[���   ;��n����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M��B$��;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P����Q�B`�Ѓ�(;��^��_^[���   ;��N����]�$ �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B�H,�у�;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B���   �у�;��[��_^[���   ;��K����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B�H(�у�;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H���   �҃�;��X��_^[���   ;��H����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��X  �у�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M���x  ��;��[��_^[���   ;��K����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�H�у�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��H  �у�;��[��_^[���   ;��K����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H��D  �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EPj�����Q�M��B��;��`���E�_^[���   ;��M����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���j �EP����Q�M��B��;������E�_^[���   ;�������]� ������������������������������������U����   SVWQ��4����3   ������Y�M���j j�����P�M��B��;��c���E�_^[���   ;��P����]��������������������������U����   SVWQ��4����3   ������Y�M��M��7��_^[���   ;�������]������������������U����   SVWQ��4����3   ������Y�M�j j �E�P�M�]����E�_^[���   ;������]� ��������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�H�у�;��>��_^[���   ;��.����]� �������������������������������������U����   SVWQ��0����4   ������Y�M���EP�M�Q����B�H�у�;������uǅ0���   �
ǅ0���    ��0���_^[���   ;������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M����   ��;����_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M�����P��M��B��;����_^[���   ;������]���������������������������������U����   SVWQ��(����6   ������Y�M��EP�M������E�M��$���_^[���   ;��)����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BX�Ѓ�;����_^[���   ;������]�������������������������U����   SVWQ��(����6   ������Y�M��EP�M��<����E�EP�M�����_^[���   ;��E����]� ����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q������   �H`�у�;���
��_^[���   ;���
����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bt��;��b
��_^[���   ;��R
����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M��Bl��;���	��_^[���   ;���	����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�hF  �EP�MQ�M�����_^[���   ;��k	����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�h#  �EP�MQ�M��Y��_^[���   ;�������]� ����������������������������������U����   SVWQ��(����6   ������Y�M���EP����Q�M����   ��;�����E�}� u3���M�����_^[���   ;��j����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �B�Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M��E��@    �E��     �E��@    �E��@   �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q@�M����   ��;����_^[���   ;������]� ��������������������������U����   SVW��@����0   ���������H|��Q ��;��?��_^[���   ;��/����]�������������������������U����   SVW��@����0   ���������H|����;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP����Q@���   �Ѓ�;��t��_^[���   ;��d����]������������������������������U����   SVW��@����0   ���������H@��Q0��;����_^[���   ;�������]�������������������������U����   SVW��@����0   ���������H@��Q0��;����_^[���   ;������]�������������������������U����   SVW��@����0   �������j�EPj ����Q@�B4�Ѓ�;��C��_^[���   ;��3����]�����������������������������U����   SVW��@����0   �������EP�MQj ����B@�H4�у�;�����_^[���   ;�������]���������������������������U����   SVW��@����0   �������j�EPh   @����Q@�B4�Ѓ�;��`��_^[���   ;��P����]��������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVW��@����0   ������h��hE  �M�������e�����Ph��hE  �M�������I���P����H��T  �҃�;��U��_^[���   ;��E����]�����������������������������������������������U����   SVW��@����0   �������EP�MQ����B��T  �у�;�����_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ������   �M����   ��;��X��_^[���   ;��H����]� �������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M��BT��;��� ��_^[���   ;��� ����]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;��o ��_^[���   ;��_ ����]�������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��B|��;�� ��_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P@�M����   ��;�����_^[���   ;��x�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��BX��;�����_^[���   ;�������]� �������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B|�H(�у�;������E�     _^[���   ;�������]������������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B|�H�у�;������E�     _^[���   ;�������]������������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B@�H�у�;������E�     _^[���   ;�������]������������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B@�H�у�;������E�     _^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ������   �M����   ��;�����_^[���   ;��|�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M��Bt��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q@�BH�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M����   ��;��+���_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ������   �M��P��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��B$��;��4���_^[���   ;��$�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP������   �M����   ��;�����_^[���   ;�������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M��Bx��;��7���_^[���   ;��'�����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��d  �у�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;��?���_^[���   ;��/�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M��Pl��;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��Bd��;��R���_^[���   ;��B�����]� �������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��Bt��;������_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M����   ��;��l���_^[���   ;��\�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M����   ��;������_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M��B��;��x���_^[���   ;��h�����]� �������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M����   ��;�����_^[���   ;��������]������������������������������U����   SVW��4����3   ������}qF t�1�E�E��}� u�#�EP�M��_���E�P�MQ�M�����������_^[���   ;��i�����]�����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q �BH�Ѓ�;������_^[���   ;��������]�������������������������������������U����   SVWQ��4����3   ������Y�M��} u�4�} t�EP�M������ �} t�EP�M�A����E�P�M�3��_^[���   ;��T�����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��B@��;������_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M����   ��;��o���_^[���   ;��_�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��BD��;������_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M�����P@��M��B`��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q@�B�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H@�Q�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P@�M����   ��;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���E P���E�$�MQ�UR�EP�MQ������   �M����   ��;�����_^[���   ;��o�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B@�HL�у�;������_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M����   ��;��{���_^[���   ;��k�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M��P\��;������_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M��Pp��;��~���_^[���   ;��n�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��Bh��;�����_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��Pp��;�����_^[���   ;��~�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M��B ��;�����_^[���   ;��������]� �������������������������������U����   SVWQ��(����6   ������Y�M���E�P����Q@�B�Ѓ�;������E�E�#Et�E��#E�E��	�E�E�E��E�P�M�Q����B@�H�у�;��O���_^[���   ;��?�����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M���D  ��;������_^[���   ;�������]� ����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B@�H�у�;��N���_^[���   ;��>�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B@�H �у�;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVW��@����0   �������j �EP����QD��Ѓ�;�����_^[���   ;��������]��������������������������������U����   SVW��@����0   �������j h�_ ����HD��҃�;�����_^[���   ;�������]��������������������������������U����   SVW��@����0   �������EPhO  ����QD��Ѓ�;��#���_^[���   ;�������]�����������������������������U����   SVW��@����0   �������j �EP����QD��Ѓ�;�����_^[���   ;�������]��������������������������������U����   SVW��@����0   �������j h:  ����HD��҃�;��F���_^[���   ;��6�����]��������������������������������U����   SVW��@����0   �������j h�  ����HD��҃�;������_^[���   ;��������]��������������������������������U����   SVW��@����0   �������EPh'  ����QD��Ѓ�;��c���_^[���   ;��S�����]�����������������������������U����   SVW��@����0   �������EP�MQ����BD��у�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EPh2  ����QD��Ѓ�;�����_^[���   ;��s�����]�����������������������������U����   SVW��@����0   �������j h�F ����HD��҃�;�����_^[���   ;�������]��������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��%����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��%����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��%����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��%����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��%����E�     _^[���   ;�������]��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;��2���_^[���   ;��"�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;��R���_^[���   ;��B�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;������_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;��r���_^[���   ;��b�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;�����_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;��"���_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;��B���_^[���   ;��2�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;������_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;��b���_^[���   ;��R�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;������_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;�����_^[���   ;��r�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;��2���_^[���   ;��"�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;��R���_^[���   ;��B�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;������_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H$�у�;��n���_^[���   ;��^�����]� �������������������������������������U���4  SVWQ�������M   ������Y�M���E�P������Q����BX�H�у�;�������   ���}�E_^[��4  ;��������]� �����������������������������������U����   SVWQ��$����7   ������Y�M��M��~����E�    �E�    �E�Pj�M�脣����u3���E�R��P�������XZ_^[���   ;��0�����]Ð   �����   �rp �������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B$�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ������;   ������Y�M���E�P�����Q����BX��у�;��,����U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��������]� �������������������������������������������U����   SVWQ������;   ������Y�M���E�P�����Q����BX�H�у�;��{����U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��C�����]� ������������������������������������������U����   SVWQ������;   ������Y�M���E�P�����Q����BX�H�у�;�������U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;�������]� ������������������������������������������U����   SVWQ��$����7   ������Y�M��} u3��0�M��4����E�    �E�E�E�Pj�M��;�����u3���   R��P�T�����XZ_^[���   ;��������]�    \�����   h�rp �����������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HD�Q�҃�;��K���_^[���   ;��;�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H �у�;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H�у�;��N���_^[���   ;��>�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H�у�;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H�у�;��N���_^[���   ;��>�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H�у�;������_^[���   ;�������]� �������������������������������������U����   SVW��@����0   ���������H\����;��`���_^[���   ;��P�����]��������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H0�у�;������_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�HH�у�;��n���_^[���   ;��^�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H�у�;������_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�HD�у�;��n���_^[���   ;��^�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q\�B�Ѓ�;������_^[���   ;��������]����������������������������U����   SVW��@����0   �������E�Q����B\�H�у�;������E�     _^[���   ;��l�����]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H\�Q8�҃�;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q\�B4�Ѓ�;�����_^[���   ;��r�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q\�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B\�H`�у�;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q\�B�Ѓ�;��"���_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H@�у�;�����_^[���   ;�������]� �������������������������������������U���  SVWQ�������B   ������Y�M��E�P�M�O����}� |o�M��H����E�P�M�5����}� tU�E�    �	�E����E��E�;E�};�E�P�M�	����E�P�M������	�Eȃ��EȋE�;E��E�P�M��r�����봸   R��P����u���XZ_^[��  ;�������]�    ������   И����   ̘����   ʘ����   Șb a cnt level ��������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H�у�;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H\�Q�҃�;��K���_^[���   ;��;�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H<�у�;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H �у�;��N���_^[���   ;��>�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H\�Q$�҃�;������_^[���   ;�������]� ����������������������������������U����   SVWQ������?   ������Y�M�j �M�6����M������EȋE�P�M�����E�    �	�E���E�E�;E�}3�E�P�M�Qh����U�R�M��:����E�P�M������E�P�M�Ԕ���R��P�X�����XZ_^[���   ;��������]�    `�����   z�����   x�b a ��������������������������������������������������������������������U���,  SVWQ�������K   ������Y�M��}}�B  �E�E��E������E�E���EE�EȋE����EE�E��}�~�E���E�E�+E�E��1�EP�M�Q�U�R�M�������E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��Y�����}�Eԃ��EԋE��E���E�P�M�Q�U���M����;��)�����}�EP�M�Q�U�R�M��(������U��������_^[��,  ;��������]� ����������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M�蕇���E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��������}�Eԃ��EԋE��E���E�P�M�Q�U���M����;�萿����}�E�P�M�Q�U�R�M���������U��������_^[��8  ;��Z�����]� �����������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U���  SVWQ�������E   ������Y�M��} t�} t�} t�} u3��  kE E�E���E�P�MQ�U���M����;��ڽ���Eȃ}� u
�E���   ��}� }3���   �E�   �E���E��E�;E���   �E�E����EԋE�E�E�E���E�P�MQ�U���M����;��i����Eȃ}� uP�}� ~C�Eԃ��EԋE�E�E�E���E�P�MQ�U���M����;��'�����t�
��E��E�뷋E��#��}� }�Eԃ��E��	�Eԃ��E��G���3�_^[��  ;��߼����]� ������������������������������������������������������������������������������������������������������U���  SVWQ�������E   ������Y�M��} t�} t�} t�} u�E� ����3���  kE E�E���E�P�MQ�U���M����;������Eȃ}� u
�E��  ��}� }�E�     3��  �E�   �E���E��E�    �E�;E���   �E�E����EԋE�E�E�E���E�P�MQ�U���M����;�耻���Eȃ}� uS�}� ~C�Eԃ��EԋE�E�E�E���E�P�MQ�U���M����;��>�����t�
��E��E�뷋E���   ��}� }�Eԃ��E��	�Eԃ��E��D����}� ~�Eԃ��M���E�Mԉ�E�;M}F�E�M�M�M���E�P�MQ�U���M����;�贺����|h�u�8���9P�6������E�8 ~I�E����MM�M���E�P�MQ�U���M����;��c�����h�u�8���?P�������3�_^[��  ;��7�����]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��u�EP�MQ�UR�M�苪���Q�} uǅ0���   �
ǅ0���    ��0�����t�EP�MQ�UR�M��������EP�MQ�UR�M��H���_^[���   ;�������]� ��������������������������������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M��Dy���E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;�葷����}�Eԃ��EԋE��E���E�P�M�Q�U���M����;��a�����}�E�P�M�Q�U�R�M��ox�����U��������_^[��8  ;��+�����]� ������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et4�E���E�Mf�f�U�E���E�M�Uf�f��Ef�M�f���_^[��]� ������������������������������������������U����   SVW��@����0   ������E;Et�&�} t �} t�} t�EP�MQ�UR�q�����_^[���   ;�襵����]�������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�跧���EP�M���訧���EP�M���0虧���EP�M���H芧���E�_^[���   ;�������]� �������������������������������������������U���L  SVWQ�������S   ������Y�M��M��d����M����Y����M���0�N����M���H�C�������s�$����s�$����s�$������苨���M����P�Q�P�Q�P�Q�P�Q�@�A����s�$����s�$����s�$�������+����M������P�Q�P�Q�P�Q�P�Q�@�A����s�$����s�$����s�$�������ȧ���M���0���P�Q�P�Q�P�Q�P�Q�@�A����s�$����s�$����s�$������e����M���H���P�Q�P�Q�P�Q�P�Q�@�A�E�_^[��L  ;��������]�������������������������������������������������������������������������������������������������������������������������������������U���  SVWQ�������C   ������Y�M��M������M����������Pv�$������肧���E���������������P�� ����H������P������H������P���`v�$������/����E���������������P�� ����H��$����P��(����H��,����P�E��@0    �E�_^[��  ;��w�����]�����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��E� �E��E�@�E��E�@�E�_^[��]� ���������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�M�P;Quljj�M��Q�����u��   �   k� �U���U���   �� �M���M�I��   ���M���M�I��   k� �U��B�   �}jj�M�������u�k�   k� �U���U���   �� �M���M�I��   ���M���M�I��   k��U���U�R��   k� �U��B�   �E�_^[���   ;��/�����]� ��������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �EP�M������E�_^[���   ;��j�����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��M��i���_^[���   ;�蘭����]������������������U����   SVWQ��4����3   ������Y�M��EP�M�踷���E�_^[���   ;��A�����]� ������������������������U���8  SVW�������N   ������j �M��T����E�M�@8�YAX�U�E�JP�YH@�\��M�YA�U�E�JP�YH(�M�U�Q �YRX�\ʋE�YH0�X��M�U�I �YJ@�E�M�P8�YQ(�\ʋU�YJH�X��E��E�f.�s���Dz�M�҃���E�  ��s�^E��E��E�M�@�YAX�U�E�JP�YH�\��M�YA0�U�E�J�YH8�M�U�Q�YR@�\ʋE�YHH�X��M�U�IP�YJ@�E�M�P8�YQX�\ʋU�Y
�X��YE��E��E�M�@�YA(�U�E�J �YH�\��M�YAH�U�E�J �YHX�M�U�QP�YR(�\ʋE�Y�X��M�U�IP�YJ�E�M�P�YQX�\ʋU�YJ�X��YE��E��E�M�@8�YA(�U�E�J �YH@�\��M�Y�U�E�J@�YH�M�U�Q8�YR�\ʋE�YH�X��M�U�I�YJ �E�M�P�YQ(�\ʋU�YJ0�X��YE��E��E�M�@8�YAX�U�E�JP�YH@�\��YE��E��E�M�@P�YA(�U�E�J �YHX�\��YE��E��E�M�@ �YA@�U�E�J8�YH(�\��YE��EċE�M�@@�YAH�U�E�JX�YH0�\��YE��E̋E�M�@X�YA�U�E�J(�YHH�\��YE��EԋE�M�@(�YA0�U�E�J@�YH�\��YE��E܋E�M�@0�YAP�U�E�JH�YH8�\��YE��E�E�M�@H�YA �U�E�J�YHP�\��YE��E�E�M�@�YA8�U�E�J0�YH �\��YE��E��   �u��}�ER��P����s���XZ_^[��8  ;�觨����]�   ������`   ��mi ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��0����4   ������E�M� �Y�U�E�J�YH�X��M�U�I�YJ�X����$�/������]��E�f.�s���Dz����s�$�M�1����E�[��s�^E��E�E�@�YE���$�M�A�YE���$�U��YE���$�M裚���E_^[���   ;��a�����]���������������������������������������������������������������������������U����   SVW��@����0   ������E�@�YE���$�M�A�YE���$�U��YE���$�M�ޙ���E_^[���   ;�蜥����]��������������������������������������U����   SVW��@����0   ������E�M�@(�Y�U�XB�E�M�H@�YI�X��U�E�JX�YH�X����$�M�U�A �Y�E�X@�M�U�I8�YJ�X��E�M�HP�YI�X����$�U�E�B�Y �M�X�U�E�J0�YH�X��M�U�IH�YJ�X����$�M記���E_^[���   ;��f�����]��������������������������������������������������������������������������������U����   SVW��@����0   ������E�M�@�\A���$�U�E�B�\@���$�M�U��\���$�M�֗���E_^[���   ;�蔣����]����������������������������������������������U����   SVW��@����0   ������E�M�@�XA���$�U�E�B�X@���$�M�U��X���$�M�&����E_^[���   ;�������]����������������������������������������������U����   SVW��@����0   ������E�M� �YA�U�E�J�Y�\����$�M�U�A�Y�E�M��YI�\����$�U�E�B�Y@�M�U�I�YJ�\����$�M�<����E_^[���   ;��������]����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M� �X�U���E��M�@�XA�U��B�E��M�@�XA�U��B�E�_^[��]� ��������������������������������������������U����   SVW��@����0   ��������E�$�ܨ����_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M��E��x0 ��   �E��M� f/v�E��M�� �E��M�@f/Av�E��M�A�@�E��M�@f/Av�E��M�A�@�E�M�� f/Av�E��M��@�E�M��@f/A v�E��M�A�@ �E�M��@f/A(v�E��M�A�@(�`�E����M���Q�P�Q�P�Q�P�Q�P�I�H�U����E��
��J�H�J�H�J�H�J�H�R�P�E��@0   _^[��]� �����������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�虈���} ��   ��h�u�<���P�M��Q����B���   �у�;�蜞���U���E��8 u3��r�} tQ��h�u�<���
P�M��Q����B���   �у�;��S����U��B�E��x u�E�P�k����3���E��M�H�E��M�H�   �3�_^[���   ;��	�����]� ����������������������������������������������������������������U����   SVW��4����3   ������j�+  ���E��}� u3���E���H��;��}���_^[���   ;��m�����]�����������������������U����   SVWQ��(����6   ������Y�M�h�   �  ���E�}� t�E샸�    u3����EP�U�M����   ��;�����_^[���   ;��ߜ����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �  ���E�}� t�E샸�    u����/��EP�MQ�UR�EP�MQ�UR�E�M����   ��;��:���_^[���   ;��*�����]� �������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S  ���E�}� t�E샸�    u����/��EP�MQ�UR�EP�MQ�UR�E�M����   ��;��z���_^[���   ;��j�����]� �������������������������������������������������U���4  SVWQ�������  ������Y�M���s�E��E�    j �M��U���j �M��K���j ��p����>����E��H�U�<�}���x  �} ��  ��P����\q��j ��0��������   k� �U��kM��U��A�E��Q�U��A�E��Q�U��A�EčE�P�   �� �U��kMQ������R�l�������0����P��4����H��8����P��<����H��@����P��D����E�   �	�E܃��Eܸ   k� �U��B�U�;��   �E�P�M���E�k�MQ�����R�-l������M��P�U��H�M��P�U��H�M��P�U��E�P��0���Q��(���R�m�����P��P��������E���0����M���4����U���8����E���<����M���@����U���D����6�������s�$��H���聎���E��H������L����P��P����H��T����P��X����H��\����P��P���P��h���Q�k�����U��H��
�H�J�H�J�H�J�H�J�@�B����P����$��[����ݝ��������������X����$��������[����ݝ����������f/������&  ����P����$�[����ݝ��������������`����$�������a[����ݝ����������f/�������   �E��HP����s�$����s�$����s�$�������ԋ��P������Q�������U����
�H�J�H�J�H�J�H�J�@�B�E��P�M��HQ������R�:������M��0���P�Q�P�Q�P�Q�P�Q�@�A��  ����X����$�iZ����ݝ��������������`����$�������;Z����ݝ����������f/�������   ����s�$����s�$����s�$������赊��P�E��HP�����Q�Y������U����
�H�J�H�J�H�J�H�J�@�B�E��P�M��HQ��(���R�������M��0���P�Q�P�Q�P�Q�P�Q�@�A�   ����s�$����s�$����s�$��H�������P�E��HP��h���Q蕋�����U��0��
�H�J�H�J�H�J�H�J�@�B�E��HP�M��0Q������R�P������M�����P�Q�P�Q�P�Q�P�Q�@�A�EP������Q������   ���}��E�    �	�E܃��E܋E�;E}�E��H�U܋E���E��ۋE���U�k�EP�MQ�����R�~�������M��P�U��H�M��P�U��H�M��P�UċE���U�kD�EP�MQ��0���R�7�������M��P�U��H�M��P�U��H�M��P�U��E�    �	�E܃��E܋E��H�U�E�;���   �E܃��M��I�u��<�UЋE��k�UR�EP��P���Q跑�������p����H��t����P��x����H��|����P�U��@�E���p���P�M�Q�U�R�  ��ݝ�����������XE��E�E��E��M��M��U��U��E��E��M��M��U��Uċ�p����E���t����M���x����U���|����E��M��M��U��U�������E�R��P�������XZ_^[��4  ;��,�����]� �I    �����   a�����   ^�p���   [�P���   Y�0���   T�prev n v3 v2 v1 ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��8����2   ������E�M�@�\A�U�Y�E�M�H�\I�U�Y
�X��E�M�H�\I�U�Y
�X���8���݅8���_^[��]���������������������������������U����  SVWQ��<����q   ������Y�M��M��f���E�    �	�Ẽ��E̋E��M�;H�	  �E���U̍��m����u�ҋE���U̍��_����E�E��E��M��P;Qud�E�kMQ�U�kBEP��@���Q��a����P�U�kEP�M�kQUR��`���P�a����P������Q������P�M��~���c�E�kMQ�U�kBEP������Q�oa����P�U�kBEP�M�kQUR������P�Ia����P������Q趄����P�M��3~��������E�P�MQ��`�����ER��P����V���XZ_^[���  ;�芎����]� �   ������   ��v ����������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j �f   ���E�}� t	�E�x  u3����EP�U�M��B ��;�訍��_^[���   ;�蘍����]� �������������������������������U����   SVW��@����0   ������h��EPh_� �s����_^[���   ;��/�����]�������������������������U����   SVWQ��(����6   ������Y�M�j<�v������E�}� t	�E�x< u���EP�U�M��B<��;�躌��_^[���   ;�誌����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�j8��������E�}� t	�E�x8 u3����E�M��P8��;��,���_^[���   ;�������]��������������������������������������U����   SVWQ��(����6   ������Y�M�jx�V������E�}� t	�E�xx u3����EP�MQ�U�M��Bx��;�蔋��_^[���   ;�脋����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��M���t���} �{  �} �q  ��h�u�D���P�M��Q����B���  �у�;������U���E��8 u3��0  �} ta�} t[��h�u�D���
P�M��Q����B���  �у�;�萊���U��B�E��x u�M��:t��3���   �E��M�H�Y�E��@   ��h�u�D���P�M��Q��R����H���  �҃�;��)����M��A�E��x u�M���s��3��p�E��M�H�E��Q�U��B��P�M��R�EP�]�����} t&�E��HQ�U��B��P�M��QR�EP�\]������   k� �U��B�U��   _^[���   ;�莉����]� ���������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��r���} �.  �E�8 �"  �E�x �  ��h�u�@���P�M�Q��R����H���  �҃�;�葈���M���E��8 u3���   �E�x tX�E�x tO��h�u�@���
P�M�Q��R����H���  �҃�;��7����M��A�E��x u�M���q��3��q�E��M�Q�P�E��M�Q�P�E��Q�U��B��P�M��R�E�Q�[�����E��x t'�E��HQ�U��B��P�M��QR�E�HQ�S[�����   _^[���   ;�蛇����]� ��������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�U�M��B��;��؆��_^[���   ;��Ȇ����]� �������������������������������U����   SVWQ��(����6   ������Y�M�jp�������E�}� t	�E�xp u3����EP�MQ�U�M��Bp��;��D���_^[���   ;��4�����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jT�f������E�}� t	�E�xT u���E�M��PT��;�讅��_^[���   ;�螅����]����������������������������������������U����   SVWQ��4����3   ������Y�M��E����   @t�����E�� %���3ҹ   ���_^[��]��������������������������������U����   SVWQ��(����6   ������Y�M�j4�f������E�}� t	�E�x4 u������EP�MQ�U�M��B4��;�裄��_^[���   ;�蓄����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M��} |�E��8 u����<�E�    �	�E���E�E��M�;H}�E���U���T��;Eu�E���Ѓ��_^[���   ;�������]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��E�P�Q�����E���P��P�����E��@    �E��@    _^[���   ;��Q�����]���������������������������U����   SVW��(����6   ������E�8 u�>j�������E��}� u�)�E��M��E�P�M��Q�҃�;��ւ���E�     R��P����x���XZ_^[���   ;�謂����]Ð   ������   ��i ����������������������������������������������U����   SVWQ��(����6   ������Y�M�j\��������E�}� t	�E�x\ u���E�M��P\��;�����_^[���   ;��������]����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �3������E�}� t�E샸�    u���EP�U�M����   ��;��q���_^[���   ;��a�����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�jh�������E�}� t	�E�xh u�(��EP�MQ�UR�EP�MQ�U�M��Bh��;��ʀ��_^[���   ;�躀����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�j(��������E�}� t	�E�x( u3����E�M��P(��;��<���_^[���   ;��,�����]��������������������������������������U����   SVWQ��(����6   ������Y�M�jP�f������E�}� t	�E�xP u3����E�M��PP��;����_^[���   ;������]��������������������������������������U����   SVWQ��$����7   ������Y�M��M��KO����E�E�M��vO����$�����$�������$�����$���w}��$����$����E� ����E� ����\�E�M���E�M�Q��E�E�M�Q��E�M�Q��-�E�M�Q��E�M�Q���E�M�Q��E�M��_^[���   ;��~����]� �I '�;�R�j�������������������������������������������������������������������������������U����   SVWQ������9   ������Y�M��E� �E�    �	�E����E��E��M�;H}3�E���U�����M��;Eu�]�E���U���������؈]���E���_^[���   ;��}����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�j$��������E�}� t	�E�x$ u2����EP�U�M��B$��;��}��_^[���   ;���|����]� �������������������������������U����   SVWQ��(����6   ������Y�M�jL�6������E�}� t	�E�xL u3����E�M��PL��;��||��_^[���   ;��l|����]��������������������������������������U���L  SVWQ�������S   ������Y�M��E��x0 ��   ���@v�$�E���P�M�Q������R������P������P�b������M���P�Q�P�Q�P�Q�P�Q�@�A�EP�M���Q������R�N�����M���P�Q�P�Q�P�Q�P�Q�@�A�{����s�$������p���E������������P�� ����H��$����P��(����H��,����P�E�M���P�Q�P�Q�P�Q�P�Q�@�A_^[��L  ;���z����]� �����������������������������������������������������������������������������������������������U���$  SVWQ�������I   ������Y�M��M��TV���E�    �	�E����E��E��M�;H��   �E���U����W����u�ҋE���U����J����E�E��E�kMQ�M��IY���E�kHMQ�M��6Y���E�kHMQ�M��#Y���E��M��P;Qt�E�kHMQ�M��Y���[����EP�MQ�M��_<��R��P����E���XZ_^[��$  ;��yy����]�    ������8   ��mm �������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j,�v������E�}� t	�E�x, u3����E�M��P,��;��x��_^[���   ;��x����]��������������������������������������U����   SVWQ������9   ������Y�M��E�    �E�    �	�E����E��E��M�;H} �E���U����kH�����t	�E���E��̋E�_^[���   ;��	x����]�����������������������������������U����   SVWQ������9   ������Y�M��E�    �E�    �	�E����E��E��M�;H}�E���U�����T����t	�E���E��͋E�_^[���   ;��jw����]������������������������������������U����   SVWQ������9   ������Y�M��E�    �E��x|�E��8 u3��?�E�    �	�E����E��E��M�;H}�E���U����E����t	�E���E��͋E�_^[���   ;��v����]�����������������������������������������������U����   SVWQ��(����6   ������Y�M��E�E��	�E���E�E��M�;H}!�E���U���pD����t�E�+E����˃��_^[���   ;��v����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�jX�F������E�}� t	�E�xX u���E�M��PX��;��u��_^[���   ;��~u����]����������������������������������������U����   SVWQ��4����3   ������Y�M��E�� %    _^[��]�����������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3����EP�MQ�U�M����   ��;��t��_^[���   ;��t����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�j��������E�}� t	�E�x u3�� ��EP�MQ�UR�E�M��P��;�� t��_^[���   ;���s����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    _^[��]��������������������������������U����   SVWQ��(����6   ������Y�M�jl�������E�}� t	�E�xl u3�� ��EP�MQ�UR�E�M��Pl��;���r��_^[���   ;���r����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�jt�������E�}� t	�E�xt u3����EP�MQ�U�M��Bt��;��Tr��_^[���   ;��Dr����]� �������������������������������������������U����   SVWQ������9   ������Y�M��M���A���E�M��B���E��E;E�t	�}���u�E;E�t	�}���u�^�}���t�E�E��}���t�E�E�}��t�E�M����E����   �ыE����E���   @�M����   �M��_^[���   ;��Hq����]� ���������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j`�f������E�}� t	�E�x` u3����EP�MQ�U�M��B`��;��p��_^[���   ;��p����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jD��������E�}� t	�E�xD u3����EP�U�M��BD��;��p��_^[���   ;���o����]� �������������������������������U����   SVWQ��(����6   ������Y�M�j0�6������E�}� t	�E�x0 u3����EP�U�M��B0��;��xo��_^[���   ;��ho����]� �������������������������������U����   SVWQ��(����6   ������Y�M�jH�������E�}� t	�E�xH u���EP�U�M��BH��;���n��_^[���   ;���n����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��Gn��_^[���   ;��7n����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3����EP�MQ�U�M����   ��;��m��_^[���   ;��m����]� ����������������������������������U����   SVW��@����0   ��������E�$��+ ��_^[���   ;�� m����]��������������������������U����   SVWQ��(����6   ������Y�M��M��=���E�}��u3��
�   �M���_^[���   ;��l����]���������������������������U����   SVWQ��(����6   ������Y�M�jd��������E�}� t	�E�xd u3����EP�MQ�U�M��Bd��;��4l��_^[���   ;��$l����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j�V������E�}� t	�E�x u3����EP�U�M��B��;��k��_^[���   ;��k����]� �������������������������������U����   SVWQ��(����6   ������Y�M�j@��������E�}� t	�E�x@ u���EP�U�M��B@��;��
k��_^[���   ;���j����]� ���������������������������������U����   SVWQ������<   ������Y�M��E�    �	�E���E�E��M�;H}�E���U��%����M���M�����E�    �	�E���E�E��M�;H}{�E���U��%   �ud�E���U���::���EԋE���E��	�E����E��E��M�;H}2�E���U����:��;E�u�E���U���   ��M���M�����q���_^[���   ;���i����]������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j|��������E�}� t	�E�x| u3����EP�U�M��B|��;��(i��_^[���   ;��i����]� �������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S������E�}� t�E샸�    u3��'��EP�MQ�UR�EP�U�M����   ��;��h��_^[���   ;��sh����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�U�M��B��;���g��_^[���   ;���g����]� �������������������������������U����   SVW��(����6   ������} t�E�8 t�E� �Pj�EP��{�����E��}� u3��5�M��|/���E�}� u3�� �} t�E�M��E�M;H~3���E�_^[���   ;�� g����]������������������������������������������U����   SVW��@����0   ������E�M��E�M�H�EPj�MQ�n����_^[���   ;��f����]����������������������������U����   SVW��@����0   ������   _^[��]�����������������������U����   SVW��4����3   ������E��M��E�M���E�M��_^[��]������������������U����   SVWQ��4����3   ������Y�M��M��VP���E�� �v�E��M�H�E�_^[���   ;��e����]� ��������������������������U����   SVWQ��4����3   ������Y�M��E�� |v�M����m���M����m���E��@    �M��V���E�_^[���   ;��e����]��������������������������������������U����   SVWQ��4����3   ������Y�M��E�� pv�E��@    �E��@    �E�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��E�� �v�M��:%��_^[���   ;��Od����]�������������������������U����   SVWQ��4����3   ������Y�M��E�� |v�M��j���M����p���M����p��_^[���   ;���c����]�����������������������������������U����   SVWQ��4����3   ������Y�M��E�� pv�M��_=��_^[���   ;��oc����]�������������������������U����   SVWQ��4����3   ������Y�M��M��T2���E��t�E�P��v�����E�_^[���   ;��c����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��N���E��t�E�P�v�����E�_^[���   ;��b����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��nn���E��t�E�P�v�����E�_^[���   ;��!b����]� ������������������������U����   SVWQ��4����3   ������Y�M��E��M��P;Qu�M��Y����u3��&�E��H�U��B�U���E��H���U��J�   _^[���   ;��a����]� �����������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E����M�A�E�M��Q�P�E��H�U�Q�E��M�H_^[��]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��@    �E����M��A�E����M��A�E��@    _^[��]���������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��B�Ѓ�;��4`��_^[���   ;��$`����]� ���������������������������U����   SVWQ��(����6   ������Y�M��M� ���E�M��Q�P�E�M��Q�P�E�    �	�E���E�E��M�;H}�E��H�U��P�M�yt����u3���͸   _^[���   ;��o_����]� ��������������������������������������U����   SVWQ������9   ������Y�M��E��x u�E��H�M��%�E��x t�E��H�U�J�M���E��H��M��}� u3��]��h�v�H���P�M���Q�U��BP����Q��  �Ѓ�;��^���E�}� u3���E��M�H�E��M��H�   _^[���   ;��p^����]����������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�    �	�E���E�E��M�;H}�E��H�U��;Eu�E���ԃ��_^[��]� ����������������������������U���   SVWQ�� ����@   ������Y�M��M��Se���E��}� tm�M��#>���E�}� tM�E��������������������� t%��j��������������;��3]���� ����
ǅ ���    �E�    �E�E�덋M��N��_^[��   ;���\����]����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E���P�*�����E��@    �E��@    �M��A    _^[���   ;��c\����]�����������������������������U����   SVWQ������9   ������Y�M��E�    �M���c���E���M��<���E��}� t�E���E���E�_^[���   ;���[����]���������������������������������������U����   SVWQ��0����4   ������Y�M��E����M�9At�U��B��0����
ǅ0���    ��0���_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H}�E��H�U���3�_^[��]� �������������������U����   SVWQ������<   ������Y�M��E�    �M��|b���E��}� tZ�E쉅����M������U���U싅���;����uǅ���   �
ǅ���    ����� t�E���M���:���E��3�_^[���   ;��<Z����]� ���������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t�M��Q�z t�E��H��0����
ǅ0���    ��0���_^[��]������������������������������������U����   SVWQ��(����6   ������Y�M��E��M;H~	�E��H�M�} }�E    �E��M��P;Qu�M��Q����u3��Z�E��H�M��	�E���E�E�;E~�E��H�U��B�U�u�L�����ԋE��H�U�E���E��H���U��J�   _^[���   ;��X����]� ��������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E�M��Q�P�E����M�A�E��H�U�Q�E��M�H_^[��]� ���������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E��M�Q�P�E�M��H�E��M�H�E��H�U��Q_^[��]� ������������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E��M�Q�P�E�M��H�E��M�H�E��H�U��Q_^[��]� ������������������������������������U����   SVWQ��(����6   ������Y�M��E;E}	�E���E�} |$�E��M;H}�} |�E��M;H}�E;Eu�/�E��H�U���E�EP�M��Zj����t�EP�M�Q�M���>��_^[���   ;��TV����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M��E��H��Q�M���;���E�}� t�E��H��Q�M��i���E�_^[���   ;���U����]��������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|3��E�E��H���U��J�	�E���E�E��M;H}�E��H�U��B�U�u�L����Ѹ   _^[��]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�����P�M��h��_^[���   ;��T����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��x t;�E��x t2�E��H�U��B�A�E��H�U��B�A�E��@    �M��A    _^[��]�����������������������������������U����   SVWQ������9   ������Y�M��M��[���E��}� t�M��c4���E�M��-���E�E���_^[���   ;��S����]������������������������������U����   SVWQ��4����3   ������Y�M��E��@    _^[��]�����������������������������U����   SVWQ��$����7   ������Y�M��EP�M���6��j�E��HQ�U��BP�MQ�M��\��R��P���f��XZ_^[���   ;��R����]� ��   �����   �sort �����������������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|3���E��H�U�E���   _^[��]� ���������������������������U����   SVWQ��4����3   ������Y�M��E��M;H}�EP�MQ�M��	O���#�E��H;M}j �M��f����EP�M��f��_^[���   ;��Q����]� ���������������������������������������U����   SVWQ��$����7   ������Y�M��EP�M��
5��j�E��HQ�U��BP�M��G��R��P�@��d��XZ_^[���   ;���P����]� ��   H����   Tsort ���������������������������������������U����   SVWQ��4����3   ������Y�M��} |$�E��M;H}�} |�E��M;H}�E;Eu�"�E��H�U��P�M��Q�E��Q�h����_^[���   ;��2P����]� �����������������������������������������U����   SVW��@����0   ������h��EPh�f �5����_^[���   ;��O����]�������������������������U����   SVW��4����3   ������j�{������E��}� t	�E��x u3����EP�MQ�U��B�Ѓ�;��IO��_^[���   ;��9O����]�����������������������������������U����   SVW��4����3   ������j��������E��}� t	�E��x u����0��E P�MQ�UR�EP�MQ�UR�EP�M��Q�҃�;��N��_^[���   ;��N����]����������������������������������������������U����   SVW������<   ������j�;������E��}� t	�E��x uǅ��������M�x��������E�E8P�M4Q�U0R�E,P�M(Q���̍UR�W���EP�M��Q�҃�4�� ����M�1���� ���_^[���   ;��M����]����������������������������������������������������U����   SVW��4����3   ������j�[������E��}� t	�E��x u3����EP�M��Q�҃�;��-M��_^[���   ;��M����]���������������������������������������U����M��L��   ��Au,�E�    �	�U����U��}�}kE��P�U�����݋E���]��������������������U��Q�M��E��M��U��: uj��������E��8}�M�k���R�uU�����E���]� �����������������������U��Q�M��E��     �M��9 uj�{������   k� �P�U�����E���]��������������������������������U����M��L������Iy,�E�    �	�U����U��}�}kE��P�K?�����݋�]�������������������������U��Q�M��E��8 uj�J������M��9}�U�k�P�~9������]����������������������U��Q�L��   ��Au,�E�    �	�U����U��}�}kE��P�HS�����݋�]����������������������������U��Q�L������Iy,�E�    �	�U����U��}�}kE��P�@>�����݋�]������������������������������U��   k� ���Q�kS����]���������������������U��} uj�������E���M��Uk�P�!S����]���������������������������U��} uj�:������E��k����Q��R����]������������������U��Ek���Q��7����]�������U��} uj�3H������E��k����Q�7����]������������������U�����]�������U��EP�MQ�UR�p ����]��������U��EPhpjj �MQ�URj�c������u�]�������������������������U��} u�EP�MQhq�	 ����]�����������������U��Q�M��E���]�������������������U��Q�M��EP�M��?Q���M��,|�E���]� �����������U����M��E�8|j�E�P�M��JQ���M��,|�E���]�������������������U��Q�M��EP�M���P���M���|�E���]� �����������U��Q�M��M������E�� �|�E���]� ���������������U��Q�M��EP�M���7���M��`|�E���]� �����������U��Q�M��EP�M��P?���M��`|�E���]� �����������U��Q�M��EP�M��7���M��p|�E���]� �����������U��Q�M��EP�M���>���M��p|�E���]� �����������U��Q�M��EP�M��O���M��P|�E���]� �����������U��Q�M��EP�M��Z���M��P|�E���]� �����������U��Q�M��EP�M���6���M���|�E���]� �����������U��Q�M��EP�M��0>���M���|�E���]� �����������U��Q�M��EP�M��:,���M���|�E���]� �����������U��Q�M��EP�M������M���|�E���]� �����������U��Q�M��EP�M���+���M���|�U��E�H�J�E���]� ���������������U��Q�M��EP��W����P�M��J���M���|�U��E�B�E���]� �������������������������U��Q�M��E�� ,|�M���$����]���������������������U��Q�M��M��$����]��������������U��Q�M��M���'����]��������������U��Q�M��M��'����]��������������U��Q�M��M��[$����]��������������U��Q�M��M��e'����]��������������U��Q�M��M������]��������������U��Q�M��M������]��������������U��]������������U��Q�M��M��2���E��t�M�Q��W�����E���]� ��������������������U��Q�M��M��K���E��t�M�Q�W�����E���]� ��������������������U��Q�M��M���Q���E��t�M�Q�`W�����E���]� ��������������������U��Q�M��M��W	���E��t�M�Q� W�����E���]� ��������������������U��Q�M��M���%���E��t�M�Q��V�����E���]� ��������������������U��Q�M��M��5���E��t�M�Q�V�����E���]� ��������������������U��Q�M��M��t!���E��t�M�Q�`V�����E���]� ��������������������U��Q�M��M��EB���E��t�M�Q� V�����E���]� ��������������������U��Q�E�E��}�ws�M��$����|�g�H}�`��}�Y�0~�R��~�K��~�D�@�=���6���/����(���!����� ���Ђ���������]�*18?FMT[bipw~����������������������������������������������������������U����M�����h�P�E�P�x9����]�����������������U���j �M��h��hR�E�P�F9����]���������������U����EP�M����h�P�M�Q�9����]�������������U����EP�M��*��h@Q�M�Q��8����]�������������U����EP�M��9��h�Q�M�Q�8����]�������������U����EP�M��hI��h�Q�M�Q�8����]�������������U����EP�M��o:��h\R�M�Q�T8����]�������������U����EP�M����h\O�M�Q�$8����]�������������U��Q�M���|��]�����������������U����*���E�h�   h��jjh   �H�����E�}� t h   ���P�E�P�������E�   �����E��E�    ����   �� ��U��}� t�E�P�3�����E��M�U���E�A�U��Q�E��A�E��]�������������������������������������������������������U���$�} u����   ���U��)���E���E�H�M��U��E܃}� u�}A|�}Z	�M�� �M�E�  �}   s:�} u�UR�5������u�E�i  ��E�H�U�Q��u�E�M  �} u"�R���M�����   ���P% �  �E��4�M�����   �U�B�H�� �  t	�E�   ��E�    �U�U�}� tN�E��%�   �   k� �D��   �� �M�L��   ��U�}�s��A���E��D� �E�   �2�   k� �E�D��E�   �}�s��xA���M��D� �E�   j�U�Rj�E�P�M�Q�U�Rh   �E�Pj �Z;����$�E�}� u�E�6�}�u�   k� �D��!��   �� �D��   k� �L������]���������������������������������������������������������������������������������������������������������������������������������U���$�} u� ���   ���U��9'���E���E�H�M��U��E܃}� u�}a|�}z	�M�� �M�E�  �}   s:�} u�UR�z:������u�E�i  ��E�H�U�Q��u�E�M  �} u"�� ���M�����   ���P% �  �E��4�M�����   �U�B�H�� �  t	�E�   ��E�    �U�U�}� tN�E��%�   �   k� �D��   �� �M�L��   ��U�}�s��<?���E��D� �E�   �2�   k� �E�D��E�   �}�s��?���M��D� �E�   j�U�Rj�E�P�M�Q�U�Rh   �E�Pj ��8����$�E�}� u�E�6�}�u�   k� �D��!��   �� �D��   k� �L������]���������������������������������������������������������������������������������������������������������������������������������U��} tj �M�!���EP�LD����]����������������U��Q�M��E��     �M��A �UR�M��b���E���]� ��������������������U��Q�M��E��M��U��E�B�E���]� ���������������U��j�h��d�    PQ���3�P�E�d�    �M�j�M��g���E�    �E�� ��M��A    �U��E�H�J�U��E�H�J�U��E�H�J�M���-��P�M�������E��UR�E�P��#�����E������E��M�d�    Y��]� ������������������������������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M�j�M��w���E�    �E�� ��M��A    �U��B    �E��@    �M��U�Qh���M�������E������E��M�d�    Y��]� ����������������������������������������������U��Q�M��E��M��E���]� ��������U��Q�M��E���]� ����������������U��Q�M��E��H�U���J�P��P�~������]����������U����M��=�� t!����E��M������E�P������֋�]��������������������������U��Q�M��E�� ��M�Q�n&�����M����8���M������]��������������U��EP�3����]����������������U����M��E��;Mtv�M�����} th�U�U��E����t�U����U���E����E��M�+M�M�h-  h�j�U�R�k������M���U��: t�E�P�MQ�U��P������E���]� ����������������������������������������������U��Q�M��M��Y$���E��t�M�Q�PI�����E���]� ��������������������U��Q�M��M��A���E��t�M�Q��	�����E���]� ��������������������U����M��E��8 t
�M���U��	�E����E��E���]����������������������U����M��E��8 u	�E�   ��E�    �E���]�������������������������U��j�h�d�    P�����3�P�E�d�    �.���E�j8h���E�Pj�^H�����E��E�    �}� t�MQ���R�M�����E���E�    �E�E��E������M����M�d�    Y��]�������������������������������������������U�졤�]�������U��j�hZ�d�    P�����3�P�E�d�    �E�    j �M��R���E�    ��9���E��}� ��   j �(�����E��E�P������M��A?   h ��M����3���U������������B��h��j�m�����E��E��}� t���Q�M���A���E���E�    �U�U��E� �E��t�M���M��B���E������M���/���E��M�d�    Y��]�����������������������������������������������������������������������������U��j�h��d�    P�����3�P�E�d�    j �M������E�    �E�H�M��}� vB�U����U��E�H�U��<� t(�E�H�U����M�Q�M�� ���P��P�L����븋E�HQ�u<�����E������M���.���M�d�    Y��]�������������������������������������������������������������U���j j ��/�����E��}� u	�E��a��E��E��M�Q�M��$�,���} t�URj �/�����E�} u	�E�����E�E�M�Q�M��,������]�����������������������������������������U��M��$�.������u�M��$�1��Pj � /����]��������������������U��j�h��d�    P�����3�P�E�d�    �*���E�h�   h���E�Pj ������E��E�    �}� t�MQ�M��a3���E���E�    �U�U��E������E�M�d�    Y��]�������������������������������������U��j�h+�d�    P�����3�P�E�d�    �j)���E�h�   h���E�Pj �������E��E�    �}� t�MQ�M������E���E�    �U�U��E������E�M�d�    Y��]������������������������������������U�������u���h�1�x%�����M���]��������������������U��j �/ �������]�������������U��Q�E�    j � ����j�r
����P�M�=���E����E��E��]�������������������������U��Q�E��M��}� t�U���M��P��P��������]���������������������U��Qj �M������h���x��������    �M��+����]����������������U��Q�EP�MQ�U�P�MQ�c������E��}� u������E���]��������������U��E�Q�UR������]����������U��EP�MQ�UR�EP�A����]��������������������U��EP�MQ�UR�EP������]��������������������U��8�]�������U��Q�   k� �����M��	�U����U��E��x t�M��;Uu�E��@���3���]������������������������������U��Q�   k� ��@��M��	�U����U��E��x t�M��;Uu�E��@���3���]������������������������������U��} t�EP�7����]����������U��} t�EP��6����]����������U���j�M�������E�@    �M�Q���U��E�M��H�}�s&�U�B�<��� t�M�Q����;Eu�뿋M�Q�E�����M�Q�� ��M�Q�� ��M��(����]������������������������������������������������U����M��E��H,�M���U���E��}� t�M��QR�E�P�MQ�U��B�Ѓ��֋�]� ����������������������������U��Q�E�x v*�M�Q�� �,�E��M�Q�E��� ��M���~��M�]���U�B0P��������]�������������������������������U����M�j �M�������E��H(�M���U��U��}� t�E���M��U�R�������ދE��@(    �M��Q,�U���E�E�}� t�M��U�E�P�������ދM��A,    ��]��������������������������������������������U����E�    �E���E��M��   �M�U��@t	�E���E�M��t	�U���U�E%;����E�E�    �	�M����M��U��<�0� t�E���0�;Mt�ًU��<�0� u	3��   �x�}� t5�E��
t-�MQj �UR�c�����E��}� t�E�P������3��l�=�}� t�M�Q��������t3��P�!�UR�E�P�MQ������E��}� u3��-�}� tjj �U�R�5�������u�E���E�P�o����3���]�����������������������������������������������������������������������������������U����E�    �E���E��M��   �M�U��@t	�E���E�M��t	�U���U�E%;����E�E�    �	�M����M��U��<�x� t�E���x�;Mt�ًU��<�x� u	3��   �x�}� t5�E��
t-�MQj �UR�������E��}� t�E�P�M����3��l�=�}� t�M�Q�5������t3��P�!�UR�E�P�MQ�t������E��}� u3��-�}� tjj �U�R��������u�E���E�P������3���]�����������������������������������������������������������������������������������U��EP�MQ�UR�������]��������U��EP�MQ�UR��*����]��������U��EP�MQ�UR�	�����]��������U��EP�M���R�EP�6����]�����������������U��EP�M����R�EP�����]�����������������U��EP�]������������������U��j h�  �EP������]���������U��EP� ]������������������U��EP�]������������������U��Q�E�8u�F�   �U�
�M��}� u�U�E�    �%�}�u�M�   ��U�:tj�"�������]�������������������������U����M�=X�
s6�X�����M��X����X��E�P��E��}� t�U�����]���������������������U��=X� u�t���$�X����X��MQ��X����]������������������������U��]����������U��EP�M�M+��]����������������U��Q�EP�M��_��P�MQ�M��R��P�4������]�����������������������U��Q�EP�MQ�n4�����Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ������Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ�������Ѕ�u	�E�   ��E�    �E���]���������������U��} t�EP��-����]����������U��} u�EP�MQhq�Y�����]�����������������U��]������������U��E;EtE�MQ�UR�EP�8������MQ�UR�EP�$������M;Ms�UR�EPhPq�������]�������������������������������U��Q�EP�MQ�������E��U��U���]����������������U��Q�EP�M�Q�?�������P�MQ�UR�EP�MQ�������]���������������������������U��Q�EP�3�����E��M�Q�UR�EP�MQ�UR�EP�MQ�:������]���������������������U��Q�E�E��	�M����M��U����t�M���E;�t�݋E�+E��]������������������������U��j�hh�d�    P��D���3ŉE�VP�E�d�    �E�    �	�E����E��MM����t'�EE���   k� �U�;�u	�M���M��j �UR�M�������E�    �E������E�   ��Eă��EċM�F����E������E� �E�    �E�    �	�Mȃ��MȋU�;U�#  �	�EЃ��EЋMM����t�EE���   k� �U�;�t�̋M�Q�M��V������t�E�P�M��C����MЉM��   �U�UĉUЋEE���   k� �U�;�t�MM����u.�}�s�EĉE���E�   �M�Q�M�������U���EȉE��[�MQ�UR�	��������u�MM��1�M������;�t(�}�s�EĉE���E�   �M�Q�M������U����E�������Eυ�t�MQ�UR���������t��v����M��M��E������M������E��M�d�    Y^�M�3��A����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M��EPj �   k� �E��R�	������M��A�URj �   k� �U�B�Q��������U��B��]�4 ����������������������U��Q�E���]������U��E]���������U����EP�W�������E�h�  hЕ�]��P�M�Q�������E��U��U�E�E���M����M��U����U��E���E�}� v�M��U���ӋE��]����������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M�������E�    ����E�|�������E�M�Q�M����E�}� t�n�}� t�U��U��`�EP�M�Q�=��������uhDq�M������hPP�U�R����.�E��E�M�����U��U�E��M�B�ЋM�Q������U�U��E������M��V���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M������E�    ����E�������E�M�Q�M�����E�}� t�n�}� t�U��U��`�EP�M�Q��������uhDq�M�����hPP�U�R�����.�E��E�M�����U��U�E��M�B�ЋM�Q�d�����U�U��E������M�����E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M��I����E�    ����E����a����E�M�Q�M����E�}� t�n�}� t�U��U��`�EP�M�Q��������uhDq�M��^���hPP�U�R����.�E��E�M�����U��U�E��M�B�ЋM�Q�$�����U�U��E������M������E܋M�d�    Y��]��������������������������������������������������������������������������U��Q�M��E��     3ɋU�f�J�E���]�����������������U��j�h8�d�    PQ���3�P�E�d�    �M��EP�M������E�    �M��Ȗ�UR�M��V����E������E��M�d�    Y��]� ���������������������������������������U��j�hh�d�    PQ���3�P�E�d�    �M��EP�M�������E�    �M����UR�M��*����E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��e����E�    �M��L��UR�EP�M�������E������E��M�d�    Y��]� ����������������������������������U��Q�M��M�������]��������������U��Q�M��E�� Ȗ�M��e�����]���������������������U��Q�M��E�� ��M��5�����]���������������������U��Q�M��E�� L��M��#���M��������]�������������U����M��E�;EtZ�M�Q�M�5��P�U�R�M��(��P����������t%3�t!j j�M��U����U�R�M����P�M�����EP�M��s����E���]� ��������������������������������������������U����M��E��x t2�MQ�U��J����E�����E�E�P�M�Q�������Ѕ�t�E�� �E���]� �����������������������������U��Q�M��E��H;Msh�  h �h,���������M��V���E��]� ����������������������U��Q�M��E��H;Msh�  h �h,��������M�����E��]� ����������������������U��Q�M��E��H��u�M������U��: uh�  h��h ��N������E��@��]������������������������������U��Q�M��E���]�������������������U��Q�M��E��8 uh  h��hh���������M�����E���]����������������������������U��Q�M��E���]�������������������U��Q�M��EP�M��������]� �������U��Q�M��EPj�M�������]� ��������������������U��Q�M��M������E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q�_������E���]� ��������������������U��Q�M��M��Q���E��t�M�Q�������E���]� ��������������������U��Q�M��EP�MQ�U�R���������]� ���������������U��Q�M���]� ���U����E�E�M��%�U���U�E�� t�M��+�U���U�E��t�M��#�U���U�E�� .�M���M�U��*�E���E��M��t�U�E��M���M�U�� 0  �U��E��tP�}�    u�E�f�.�}� 0  u�E�A��}�   u�E�E��E�G�M��M��U��U��E�M���U���U��N�}�    u�E�f�.�}� 0  u�E�a��}�   u�E�e��E�g�E��E��M��M��U�E���M���M�U�� �E��]����������������������������������������������������������������������������������U��j�h��d�    P���   ���3ŉE�SP�E�d�    h`  hx��EP�
�����}0 v�M ���+t�E ���-u	�E�   ��E�    �U��U��M�i��% 0  = 0  tǅ|��� ��Jǅ|���$��E���;E0w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M���|���R�   k� M Q������E�f�(�f�U�������   k� � �   k� ��T��   k� �T�R�   k� M Q�m�����E���`���R�M�	�����l�����l�����\����E�    ��\���Q�������E��E�������`�������j0�M��>���E�j �U0R�M�������E�   j �M�����P�E E0P�   k� U R�M�������p���P�M�u�����d�����d�����h����E���h���R�,�����E��E���p��������E�P�M��c���E��M������E��M$�M��U�;U0u �E�E��E��M�Q�U$R�E�P�M�����c�M�M��M��U�R�E,P�M�Q�M�����U�R�E(P�M���Q�M��k���M������؋U�R�M��������E�P�M$Q�U�R�M��>��j �M������E��E����tY�U����~O�M���E�+E�;�s?�M���E�+E��M�Qj�U�R�M������   �� �M����~	�E����E�뜍M��q����E0�M�������t�����x�����x��� |(	��t��� v�M����;E0v�M����+E0�E���E�    �M��M��M�@��%�  �E��}�@ty�}�   tp�U�R�EP�MQ�UR��<���P�MQ��������@�U�E�E�    �M�Qj �M��}���P�UR�EP��T���Q�UR��������P�M�U�   �}�   um�E�Pj �M��:���P�MQ�UR��,���P�MQ�L�������@�U�E�M�Q�UR�EP�MQ��D���R�EP���������P�M�U�E�    �5�E�Pj �M������P�MQ�UR��4���P�MQ���������@�U�E�M0+M�Q�U�R�M�����P�EP�MQ��L���R�EP��������P�M�Uj j �M������E�P�MQ�UR�EP�MQ�UR�M������E��M������E������M��}����E�M�d�    Y[�M�3��+�����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hd�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h  h`��M�Qj�m������E��E�    �}� t:j �M����P�M��y����E��U��U��E��E����E��M�Q�M��l����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ����E�hD  h`��M�Qj�-������E��E�    �}� t:j �M���P�M��9����E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��e���   �M�d�    Y��]��������������������������������������������������������������������������U��j�hD�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �m���E�h�   h`��M�Qj��������E��E�    �}� t<jj �M�W��P�M�������E��U��U��E��E����E��M�Q�M��C����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��#���   �M�d�    Y��]������������������������������������������������������������������������U���`���3ŉE�VW�M̍E�P�	�����   ���}��   �uЋ}�E_^�M�3�������]� ���������������������������������U��Q�M������]�����������������U��j�h��d�    P��   ���3ŉE�VP�E�d�    �M���% 0  = 0  u%�EP�MQ�UR�EP�MQ�UR�^������  ��\���P�M������l�����l�����d����E�    ��d���R�q�����E��E�������\����a����E�P�M������E�   �M�M��E� ��`���R�M�T�����h�����h�����p����E���p���Q���������x����E���`���������U�R�   k����Q�   k� �P��x��������MQ�UR�E���������t�h�M������Ⱥ   k��T�;�u�E�� +�M����M��M�<����3�M�����и   k�
�D�;�u�M��-�U����U��M�����E� �E�    �E�    j �M�������E��E����t�U������   ��E��M������MQ�UR����������te�M�$�����Q�U�R�A������E��}�
sD�}�$|�E����E��.�}� u�}� u� �M��U������M����M��U����U��x����  �M��������u�E� ��M��(����E��E��E�j j�M������E��E�    ��M������MQ�UR�������������   �M�[�����Q�U�R�x������E��}�
s~�E��}�$|�E����E��.�}� u�}� u� �M��U������M����M��U����U��E�P�M���������t%�U�R�M��������|�����|��������|����
�G�E�P�M��������t�U���t�M�������M�;�t��j j�M�������U����U�������}� u�"�E�P�M��d������~�U����U���E��E���u�}� vy�M����u�l�e�E����E�t�M��1�U�R�M������ ;�u�}� u�M��1�U�R�M������� ;�}�E���   �� �U��
��~	�M����M��y����E��M������U���t�}� u�E�� 0�M����M��UR�EP�������ȅ�tB�M�������M��\�����;�u(������   k� � �M����E����E��M������}� uj��E��M�����MQ�UR����������t'�M�����Ⱥ   k� �T�;�u�E����E�붃}� }�M��0�U����U��E����E���E��M�E����MQ�UR�1���������tI�M������Q�U�R��������E��}�
s(�}�$} �E��M������E����E��M����M���U�����  �EP�MQ��������Ѕ���  �M�8������   k��L�;�t �M�����и   k��D�;��i  �M��e�U����U��M�k����E� �E�    �EP�MQ�������Ѕ�t�h�M��������   k��L�;�u�U��+�E����E��M�����3�M�����Ⱥ   k�
�T�;�u�E�� -�M����M��M������UR�EP��������ȅ�t*�M�B����и   k� �D�;�u�E��M������M���t�U��0�E����E���E��M�y����MQ�UR�e���������tI�M�������Q�U�R��������E��}�
s(�}�} �E��M������E����E��M����M���U���u�E���u�M�M��U�� �E���t����E������M��������t����M�d�    Y^�M�3��k�����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��   ���3ŉE�VP�E�d�    ��P���P�M�������`�����`�����X����E�    ��X���R�������t����E�������P���臽���E�P��t���������E�   ��T���Q�M������\�����\�����d����E���d���P���������l����E���T����(����M�Q�   k�t�P�   k� ��t�R��l����G����E�E��E� �MQ�UR�h���������t�h�M�����Ⱥ   k��T�;�u�E�� +�M����M��M�_����3�M������и   k��D�;�u�M��-�U����U��M�*����E�� 0�M����M��U��x�E����E��E� �E�    ǅ|���    �MQ�UR����������u�M�Z����Ⱥ   k� �T�;�t�b�EP�M����P�������ȅ�tB�M� ����и   k��D�;�t�M�����Ⱥ   k��T�;�u
�M�f�����E�j �M��;�����x�����x������t��x��������   ��E��M�#����MQ�UR����������tk�M������Q�U�R�������E��}�sJ�}�$|��|�������|����.�}� u�}� u� �M��U���t���M����M��U����U��r����.  �M��R�����u�E� ���t��������E��E��E�j j�M�������E��E�    ��M�U����MQ�UR�A�����������   �M������Q�U�R��������E��}���   �E��}�$|��|�������|����.�}� u�}� u� �M��U���t���M����M��U����U��E�P�M��B������t%�U�R�M��.�����p�����p��������p����
�G�E�P�M��������t�U���t�M��������M�;�t��j j�M��0����U����U�������}� u�"�E�P�M��������~�U����U���E��E�����   �}� ��   ��x������u�{�t�E����E�t��x����1�U�R�M��U���� ;�u"�}� u"��x����1�U�R�M��3���� ;�}�E��%�   �� ��x����
��~��x�������x����_����E��M��I����U���t�}� u�E�� 0�M����M��UR�EP�=������ȅ�tE�M��������t���莸����;�u(������   k� � �M����E����E��M������}� uy��E��M������MQ�UR�����������t-�M�D����Ⱥ   k� �T�;�u��|�������|���밃�|��� }�M��0�U����U���|�������|�����E��M�h����MQ�UR�T���������tI�M�������Q�U�R��������E��}�s(�}�$} �E��M���t���E����E��M����M���U�����  �EP�MQ��������Ѕ���  �M�[������   k��L�;�t �M�?����и   k��D�;��i  �M��p�U����U��M�����E� �E�    �EP�MQ�@������Ѕ�t�h�M��������   k��L�;�u�U��+�E����E��M�7����3�M�����Ⱥ   k��T�;�u�E�� -�M����M��M�����UR�EP��������ȅ�t*�M�e����и   k� �D�;�u�E��M�������M���t�U��0�E����E���E��M�����MQ�UR����������tI�M�������Q�U�R�������E��}�s(�}�} �E��M���t���E����E��M����M���U���u�E���u�M�M��U�� �E��|����ǅh���    �E������M��������h����M�d�    Y^�M�3�������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hp�d�    P��   ���3ŉE�VP�E�d�    �EP� ������x����M�Q��x���������E�    �M��������u�E� ���x����,����E��U��U��EP��������X����M�Q�   k��P�   k� ���R��X����u����E�E��MQ�UR����������t�h�M�>����Ⱥ   k��T�;�u�E�� +�M����M��M葼���3�M�	����и   k��D�;�u�M��-�U����U��M�\����E%   �E�}   u	�E�   �F�}   uǅd���   �(�} uǅl���    �
ǅl���
   ��l�����d�����d����U��E��E��E� �E� �MQ�UR�������������   �M�J����Ⱥ   k� �T�;���   �E��M褻���EP�MQ�������Ѕ�tY�M�������   k��L�;�t�M������и   k��D�;�u!�}� t�}�u�E�   �E� �M�6�����}� u�E�   �}� t0�}�
t*�}�uǅt���   �
ǅt���   ��t�����h����
ǅh���
   ��h�����`����E�Pj�M��C����E��E�    �   k�U��\�����M覺���EP�MQ�������Ѕ���   �M������P�M�Q�"�������p�����p���;�`���sz�E���p��������E���u�M����0t�E�;�\���s�M����M��E��E��U�R�M�蕺��� ��t$�M�Q�M�聺����|�����|������|�����G�U�R�M��[���� ��t�M���t�M�D������E�;�t��j j�M������M����M�������}� u�"�U�R�M������ ��~�M����M���E� j �M��J����E��U���t�}� vy�E����u�l�e�U����U�t�E��0�M�Q�M�誹���;�u�}� u�E��0�M�Q�M�苹���;�}�E� ��   �� �M����~	�E����E��y����M���t�U���u�E�� 0�M����M���U���u�E�E��M�� �U���T����E� �M��l����E������M��]�����T����M�d�    Y^�M�3�������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M��������]�����������������U��Q�M��M���,������]�����������U��Q�M��ȕ��]�����������������U����E�E��M��%�U����U��E�� t�M��+�U����U��E��t�M��#�U����U��   k� �U�
��Lt�   k� �E��M���E����E��-�M��I�U����U��E�� 6�M����M��U��4�E����E��M��   �M�}�   u�E�o�:�}�   t�   �� �E��M���U��t�E�X��E�x�E��E��M��M��U��E���M����M��U�� �E��]��������������������������������������������������������������������������������������U����M��E��8 t,�M��	藶���E������E�U�R�E�P�_������ȅ�t�U��    �E��@��M��A ��]�����������������������U��Q�M���]� ���U��Q�M���]� ���U��j�h��d�    PQ��   ���3ŉE�SVWP�E�d�    �e��M��M�E����E��E�P�M�=����M��A    �U��B    �E��@    �E�    �M��t	�E��a�	�U��B�E��M�Q�M�������p�����p���Rj �E�P迹������x����M���x����Q�M�~����E��E�Pj �M�Q萹������|����U���|����B�M������t����M�Qj ��t���R�[������E��E��M��H��M�����j j �O����dy��E�������E������U��t.�E�Pj j.�}������M��A�U�Rj j,�g������M��A���,�   �u����U�Rj �M������M�d�    Y_^[�M�3�������]� ��������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��   ���3ŉE�P�E�d�    h�  hx��EP�������}$ v�M ���+t�E ���-u	�E�   ��E�    �U��U��M�����%   =   u@�E���;E$w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M��U�R�M������|�����|�����t����E�    ��t���Q�������E��E������M�赦��j �U$R�M��׼���E�   j �M��ѱ��P�E E$P�   k� U R�M�������E�P�M������x�����x����M��E��U�R�J������E��E��M��@����E�P�M������E�j �M��Ĳ���E��M����ty�E����~o�M�������E��U����tY�M����~O�E���U$+U�;�s?�E���U$+щU$�E�Pj�M$Q�M������   �� �E����~	�U����U�뜍M������E$�M�m����E��U��}� |%�}� v�M�Q���;E$v�M�D���+E$�E���E�    �E��E��M�����%�  �E��}�@ty�}�   tp�M�Q�UR�EP�MQ��T���R�EP�T�������P�M�U�E�    �E�Pj �M��&���P�MQ�UR��l���P�MQ�8�������@�U�E�   �}�   um�M�Qj �M�����P�UR�EP��D���Q�UR���������P�M�U�E�P�MQ�UR�EP��\���Q�UR覮������P�M�U�E�    �5�E�Pj �M��v���P�MQ�UR��L���P�MQ舧������@�U�E�M$+M�Q�U�R�M��<���P�EP�MQ��d���R�EP�N�������P�M�Uj j �M蜷���E�P�MQ�UR�EP�MQ�UR��������E��M��5����E������M��&����E�M�d�    Y�M�3��������]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hX�d�    P�����3�P�E�d�    j �M������E�    �E�(   �E�H;M��   �U���U��}�(s�E�(   h�   h��j�E���P�M�QR�n������E�}� u������E�M�H��U�B���M�A�U�B;E�s�M�Q�E�H��    �ыU��M�P�ҋE�H�U�<� t(�E�H�U���M�Q�M� ���P��P�������E�H�U�E���E������M��]����M�d�    Y��]������������������������������������������������������������������������������������U��j�h��d�    P��D���3�P�E�d�    �E;��u<h ��M��1����E�    j �MQj?�U�R�$������E������M������   j �M��B����E�   �E�x v}jhh��j�M�Q��R�П�����E�E�M�H�}� u�G����U�B�E��}� v<�M����M��U�B�M����U�E�H�U��E���}� t�M��M�B����E������M�������M�d�    Y��]��������������������������������������������������������������������������������U����E�    �} u
hTa腪���   k� �U�
��*u�   �� �U�
��u�|�} uj j �������E��e�}?u�MQj �������E��L�E�    �	�U����U��}�#�   �M�����#Et�MQ�U�R�L������΋EPj �<������E��}� uh���M��,蝮���,h���M��,����P�q�������t�M�Q�M��,�o����E��]��������������������������������������������������������������������U���j j �������E��}� u	�E��a��E��E��M�Q�M��$�����UR�EP�MQ��������]��������������������������������U��j�h8�d�    P��P���3�P�E�d�    j j �Z������   ������#Uu�   �} um�#����E�jJh���E�Pj覰�����E��E�    �}� tj �MQ�M��.����E���E�    �U�U��E������������P�E�P�M����� ��������P�MQ菿����P�M����j j �h������   ������#Uu�   �} um�o����E�jKh���E�Pj�������E��E�   �}� tj �MQ�M������E���E�    �U�U��E������|��[���P�E�P�M�X���� �|��B���P�MQ������P�M�6���j j �������   ������#Uu�   �} um�����E�jLh���E�Pj�>������E��E�   �}� tj �MQ�M�� ����E���E�    �U܉U��E��������觧��P�E�P�M褶��� ���莧��P�MQ�������P�M肶��j j ��������   ������#Uu�   �} uo�����E�jMh���E�Pj芮�����E��E�   �}� tj j �MQ�M������E���E�    �UԉU��E������������P�E�P�M����� ����ئ��P�MQ������P�M�̵��j j �������   ������#Uu�   �} um�Q����E�jOh���E�Pj�ԭ�����E��E�   �}� tj �MQ�M��W����E���E�    �ỦU��E������ ��=���P�E�P�M�:���� � ��$���P�MQ������P�M�����UR�EP�MQ�UR�&������EP�MQ�UR�EP��������MQ�UR�EP�MQ�������U�BE�M�A�M�+���P�M��蟩���E�M�d�    Y��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��E��8 t,�M��	�&����E�������E�U�R�E�P�?������ȅ�t�U��    ��E�P�K������M��A�U��B�E��@��]��������������������������������������U����E���E�M耗���M���M�} v�U�P�M�������+����ȋM�U��E�A�E]���������������������������������U����E���E�M�����} v�MQ�M�R�����������ӋU�E��M�J�E]����������������������������U��Q�M��E��8 tj�M��R�������E��     ��]���������������������U��Q�M��E��HQ�������U��BP�ѵ�����M��QR�µ������]�������������������������U����M��E�;Eu�a�M�Q�M����P�U�R�M��
���P����������t�M�yr�UR�M��Y����!j j�M������EP�E�����P�M�螠���E���]� �����������������������������������U��Q�M��@aPj �MQ�M��8�����]� ���������������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E��@��]����������������U����M��E�    �E��HQ�M�����U����U��E��]� ���������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP��������E�    �M�Q�M�����E��U��U��E�    �E�P�M�I���P�MQ�UR�E�P�M�Q蹝�����E��E������M��{����   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R��������E̍EP�MQ谻�����Ѕ�t�E ����U �
�E�;E�t�}� u	�}���  v�M ����E ��,�   k� �DЃ�-u
3�+M̉M���ỦUċE$f�M�f��U�E��M�J�E�M�d�    Y�M�3��������]�  ������������������������������������������������������������������������������������������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP��������E�    �M�Q�M�����E��U��U��E�    �E�P�M�Y���P�MQ�UR�E�P�M�Q�ɛ�����E��E������M�苒���   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R�������E̍EP�MQ��������Ѕ�t�E ����U �
�E�;E�t�}� u�}��v�M ����E ��*�   k� �DЃ�-u
3�+M̉M���ỦUċE$�Mĉ�U�E��M�J�E�M�d�    Y�M�3�������]�  �����������������������������������������������������������������������������������������������������������U��j�h�d�    P��@���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP��������E�    �M�Q�U�R�M������E��E��E��E�    �M�Q�M�e���P�UR�EP�M�Q�U�R�ՙ����P�E�P�M�Q蝶�����E��E������M�膐���UR�EP��������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3��r�����]�  �������������������������������������������������������������������������������U��j�hH�d�    P��@���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP�l������E�    �M�Q�U�R�M�}����E��E��E��E�    �M�Q�M�����P�UR�EP�M�Q�U�R�U�����P�E�P�M�Q�ѿ�����E��E������M������UR�EP�|������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3�������]�  �������������������������������������������������������������������������������U���T���3ŉE��M�h)  hx��EP�MQ�UR�EP�������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q质����P�U�R�E�P�9������]��}� t�M���QQ�E��$�+������]��UR�EP�������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3�蟯����]�  ����������������������������������������������������������������������������U���X���3ŉE��M�hA  hx��EP�MQ�UR�EP�������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q�d�����P�U�R�E�P�б�����]��}� t�M���Q���E��$�&������]��UR�EP�̳�����ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��M�����]�  ��������������������������������������������������������������������������U���X���3ŉE��M�hY  hx��EP�MQ�UR�EP�d������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q������P�U�R�E�P�˺�����]��}� t�M���Q���E��$�ų�����]��UR�EP�|������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��������]�  ��������������������������������������������������������������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�hq  hx��EP�MQ�UR�EP��������E�    �M�Q�M�����E��U��U��E�    �E�Ph   �MQ�UR�E�P�M�Q�������E��E������M�诉���   ��t"�E�P�M�Q�U�R�E�P�G�����3ɉE��M���U�R�E�P�M�Q�U�R�������E��U��E��E��M��M��UR�EP�а�����ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E��M$��U�E��M�J�E�M�d�    Y�M�3��F�����]�  ���������������������������������������������������������������������������������������������������U��j�h��d�    P��D���3ŉE�P�E�d�    �M�h   hx��EP�MQ�UR�EP�,������E�    �M�Q�U�R�M�=����E��E��E��E�    �M�Q�M����P�UR�EP�M�Q�U�R������P�E�P�M�Q蛸�����E��U��E������M��Ç���UR�EP�9������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3�詩����]�  ��������������������������������������������������������������������������������������U��j�h�d�    P��D���3ŉE�P�E�d�    �M�h  hx��EP�MQ�UR�EP�������E�    �M�Q�U�R�M譭���E��E��E��E�    �M�Q�M����P�UR�EP�M�Q�U�R腏����P�E�P�M�Q��������E��U��E������M��3����UR�EP詭�����ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3�������]�  ��������������������������������������������������������������������������������������U��j�hq�d�    P��   ���3ŉE�P�E�d�    ��L���h�  hx��EP�MQ�UR�EP������ǅx��������M����% @  �'  ��H���Q�M������\�����\�����P����E�    ��P���P��������p����E�������H���裄��j j�M��ǚ���E�   ��|���Q��p����o�����@�����@�����8����E���8���P�M��ɇ���E���|����ޕ��j �M�������M�Q��p���������d�����d�����<����E���<���P�M��|����E��M�蔕���M��y���Pj�MQ�UR��������x����E������M��d����   ǅh���    ��h���P��`���Q�M�ʪ����T�����T�����D����E�   ��D���P�M�&���P�MQ�UR�E�P��L���Q蓌����P��X���R�E�P��������l����E�������`����;����M�9�X���t��h��� u��l���w��l�����x����EP�MQ航�����Ѕ�t�E ����U �
��x��� }�E ����U �
�*��x��� tǅt���   �
ǅt���    �E$��t�����U�E��M�J�E�M�d�    Y�M�3�������]�  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��E�    �E��HQ�M�{����U����U��E��]� ���������������U���P���3ŉE��M��EP�M����Phؗ�M�Q�U�R�D�����Pj@�E�P�������P�M�Q�UR�EP�MQ�UR�EP�M�Q�+����� �E�M�3��f�����]� �����������������������������������U���P���3ŉE��M��EP�M�f���Phܗ�M�Q�U�R褂����Pj@�E�P�^�����P�M�Q�UR�EP�MQ�UR�EP�M�Q苢���� �E�M�3��Ƣ����]� �����������������������������������U���   ���3ŉE���`����M������T�����X�����X��� 0|	��T��� w%�M����%    uǅh���   ǅl���    ��M�g�����h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M�����% 0  =    �  �E�@v�E������D��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E������u��x����  s�E�5���]���E��s����Aud���t�����
��t����}� |M	��|���
rB�Й�]����u2��t����  s&�E����]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M����Pj �E�P��`���Q�����Pjl�U�R襻����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P苍����,�E�M�3��������]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE���`����M�T�����T�����X�����X��� 0|	��T��� w%�M�<���%    uǅh���   ǅl���    ��M������h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M����% 0  =    ��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E������u��x����  s�E�5���]���E��s����Aud���t�����
��t����}� |M	��|���
rB�Й�]����u2��t����  s&�E����]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M�f���PjL�E�P��`���Q��{����Pjl�U�R�^�����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P�D�����,�E�M�3�讜����]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���H���3ŉE��M��EPh�j@�M�Q�8�����P�U�R�EP�MQ�UR�EP�MQ�U�R�e����� �E�M�3�蠛����]� �����������������������������U���P���3ŉE��M��E P�MQ�M����Ph���U�R�E�P��z����Pj@�M�Q蚶����P�U�R�EP�MQ�UR�EP�MQ�U�R�ǚ���� �E�M�3�������]� �����������������������������������������������U���P���3ŉE��M��E P�MQ�M�����Ph��U�R�E�P�0z����Pj@�M�Q������P�U�R�EP�MQ�UR�EP�MQ�U�R������ �E�M�3��R�����]� �����������������������������������������������U��j�h��d�    P��   ���3ŉE�VP�E�d�    �M�h�  hx��EP腮�����M����% @  u4�MQ�UR�EP�MQ�UR�EP�M���M��B$�ЋE��  ��  ��p���Q�M�J����E��U���|����E�    ��|���P�������E��E�������p�����v���M��f����E�   �M��t%�U�R�M�跸���E��E�P�M��a}���M��N����#�M�Q�M�蝣���E��U�R�M��<}���M��)����M�n�����t�����x�����x��� |:	��t��� v/�M�F������M��ҋ��;�v�M�0������M�輋��+��u���E�    �E��E��M�̾��%�  ��@t6�M�Q�UR�EP�MQ��`���R�E�P�D�������P�M�U�E�    �M��X���P�M��Y���P�EP�MQ��h���R�E�P�%y������P�M�Uj j �M�s����E�P�MQ�UR�EP�MQ�U�R�������E������M��	����E�M�d�    Y^�M�3�跗����]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M��E��@��]����������������U����M��E�    �E��HQ�M�K����U����U��E��]� ���������������U����M��E��H��u�M��ʏ���U�B��u�M跏���M��9 u�U�: t�E��8 t�M�9 u	�E�    ��E�   �E���]� ����������������������������������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�P�M������P�M豔���E��]� ���������U��j�h�d�    P�����3�P�E�d�    �E�    �M��޼���E�    j �M������E�衷���E��E�M�;��   �U���M��P��P�l������E��M��U�R�K������E���M��B�ЋM��Q��?�U�}�?u�M����>���Pj �-������C�E�    �	�E���E�}�+�   �M�����#U�t�M��������P�E�P�������ƍM�Q�M诡���U����U��E� �M��W����E������M��r���E��E������M��r���M�d�    Y��]�������������������������������������������������������������������������������������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E��H;Ms�M�艦���U��@a+B;Ew�M�襚���} vo�M��QU�U�j �E�P�M���{���ȅ�tN�U��B+EP�M��ʖ��EP�M�辖��EEP��~�����MQ�UR�EP�M���n���M�Q�M��P���E���]� ����������������������������������������������U��Q�M��M��A�Q��]�������������U����M��M�������E�U��}� |,�}� v$�M��x}���E��E��M��U�R�������E���EP�������P�M���M��B�ЉE�E��]� ���������������������������������U��Q�M��E���M��B�Ћ�]���������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��EP�MQ�UR�E���M��B�Ћ�]� ����������U����M��E��H �M�P$�U��E��M�H �U�P$�E�U���]� �������������U��Q�M��M��A �Q$��]�������������U��Q�EP�E���$�m�����]��E���]��������������U��EP���E�$�gm����]�������U���8���3ŉE�VW�E�    3��EԉE؉E܉E��E�E�E�E��E�E�螗���E��
����E��cr���   ��< u	�E�   ��E�    �UȉU؃}� uQ�E�    �	�Ẽ��É}�   }6�M�Q�c������t$�U����M̃��   ���L�ȋU����L�븹   �uЋ}�E_^�M�3��	�����]�������������������������������������������������������������������������U���d���3ŉE�VW�E�x t0�M���   ~�-���� *   ����   �U�E��   �t�r�E�    �} u�M�Q艭�����   ���}��UЉU�E�Pj �M�QR�EPj�MQj �U�P��Ẽ}� t�}� t誶��� *   �����E�_^�M�3�������]����������������������������������������������������U��EP�MQ�UR�EP�������]�������������������U��]����������U��EP�M�Ý��]����������������U��Q�EP�M�����P�MQ�M��ڼ��P莊������]�����������������������U��Q�EP�M��q���P�MQ�M��d���P�ӌ������]�����������������������U��EP�M�ť��]����������������U��]����������U��Q�EP�MQ��������Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ�Œ�����Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ�z�����Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ�>������Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ�u�����Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ�5������Ѕ�u	�E�   ��E�    �E���]���������������U��Q�E�    �} u�%�}���w�E��P�V������E��}� u��x���E���]������������������U��Q�E�    �} u�%�}���w�E��P�������E��}� u�wx���E���]������������������U��Q�EP�MQ�|�����E��U�R�EP�MQ�UR�EP�MQ�������E��]������������������U��Q�EP�M�Q�t�����UR�E�P�i�����M�Q�U�R�EP�MQ�UR�EP�MQ�j������E��]��������������������������������U����M�����E���E�M;Mt�U�P�M�~����������ϋM�U��E�A�E]������������������������U��EP�MQ�UR�EP�MQ�ۂ�����E]�������������U��Q�EP�MQ�Ih�����E��U�R�EP�MQ�UR�EP�MQ�x������E��]������������������U��Q�EP�M�Q��l�����UR�E�P�Mh�����M�Q�U�R�EP�MQ�UR�EP�MQ�m������E��]��������������������������������U����M��t���E���E�M;Mt�U�P�M�u������8����ϋM�U��E�A�E]������������������������U��EP�MQ�UR�EP�MQ�ߴ�����E]�������������U��} u�EP�MQhq��{����]�����������������U��} u�EP�MQhq�{����]�����������������U��} u�EP�MQhq�{����]�����������������U��} u�EP�MQhq�Y{����]�����������������U��} u�EP�MQhq�){����]�����������������U��]������������U��]������������U��} u�EP�MQhq��z����]�����������������U��} u�EP�MQhq�z����]�����������������U��E;EtE�MQ�UR�EP�q������MQ�UR�EP�]������M;Ms�UR�EPhPq�Gz����]�������������������������������U��E;EtE�MQ�UR�EP荕�����MQ�UR�EP�y������M;Ms�UR�EPhPq��y����]�������������������������������U��E;EtE�MQ�UR�EP�4������MQ�UR�EP� ������M;Ms�UR�EPhPq�gy����]�������������������������������U��E;EtE�MQ�UR�EP�������MQ�UR�EP��������M;Ms�UR�EPhPq��x����]�������������������������������U��E;EtE�MQ�UR�EP��������MQ�UR�EP�������M;Ms�UR�EPhPq�x����]�������������������������������U��Q�EP�MQ襊�����E��U��U���]����������������U��Q�EP�MQ�m�����E��U��U���]����������������U��Q�EP�M�Q���������P�MQ�UR�EP�MQ��r������]���������������������������U��Q�EP�M�Q蒫�������P�MQ�UR�EP�MQ��}������]���������������������������U��Q�EP�M�Q�b�������P�MQ�UR�EP�MQ��������]���������������������������U��Q�EP�M�Q�l�������P�MQ�UR�EP�MQ裆������]���������������������������U��Q�EP�M�Q�,q�������P�MQ�UR�EP�MQ�rv������]���������������������������U��Q�EP�%h�����E��M�Q�UR�EP�MQ�UR�EP�MQ�+�������]���������������������U��Q�EP�Kj�����E��M�Q�UR�EP�MQ�UR�EP�MQ�v������]���������������������U��Q�E�E��	�M����M��U����t�M���E;�t�݋E�+E����]����������������������U��Q�E�E��	�M����M��U����t�M���E;�t�݋E�+E����]����������������������U��j�hH�d�    P��D���3ŉE�VP�E�d�    �E�    �	�E����E��MM����t'�EE���   k� �U�;�u	�M���M��j �UR�M��uu���E�    �E������E�   ��Eă��EċM�����E������E� �E�    �E�    �	�Mȃ��MȋU�;U�#  �	�EЃ��EЋMM����t�EE���   k� �U�;�t�̋M�Q�M���i�����t�E�P�M���i���MЉM��   �U�UĉUЋEE���   k� �U�;�t�MM����u.�}�s�EĉE���E�   �M�Q�M��ri���U���EȉE��[�MQ�UR����������u�MM��1�M�|z����;�t(�}�s�EĉE���E�   �M�Q�M��i���U����E�������Eυ�t�MQ�UR�y���������t��v����M��M��E������M��#o���E��M�d�    Y^�M�3�������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��D���3ŉE�VP�E�d�    �E�    �	�E����E��MM����t'�EE���   k� �U�;�u	�M���M��j �UR�M��r���E�    �E������E�   ��Eă��EċM荡���E������E� �E�    �E�    �	�Mȃ��MȋU�;U�#  �	�EЃ��EЋMM����t�EE���   k� �U�;�t�̋M�Q�M���f�����t�E�P�M���f���MЉM��   �U�UĉUЋEE���   k� �U�;�t�MM����u.�}�s�EĉE���E�   �M�Q�M��f���U���EȉE��[�MQ�UR�	f��������u�MM��1�M臋����;�t(�}�s�EĉE���E�   �M�Q�M��%f���U����E�������Eυ�t�MQ�UR�e��������t��v����M��M��E������M��3l���E��M�d�    Y^�M�3���|����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��D���3ŉE�VP�E�d�    �E�    �	�E����E��M��U�J��t(�M��U�J�   k� �M�;�u	�E���E��j �MQ�M��o���E�    �E������E�   ��Uă��UċM�9����E������E� �E�    �E�    �	�Eȃ��EȋM�;M�(  �	�UЃ��UЋEЋM�A��t�EЋM�A�   k� �E�;�t�ʋU�R�M��d��� ��t�M�Q�M���c���UЉU��   �E�EĉEЋMЋU�J�   k� �M�;�t�EЋM�A��u.�}�s�EĉE���E�   �M�Q�M��c���U���EȉE��\�MQ�UR����������u�MЋU�4J�M�t����;�t(�}�s�MĉM���E�   �U�R�M��.c���M����E�������Uυ�t�EP�MQ������Ѕ�t��q����E��E��E������M��<i���E��M�d�    Y^�M�3���y����]����������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��D���3ŉE�VP�E�d�    �E�    �	�E����E��M��U�J��t(�M��U�J�   k� �M�;�u	�E���E��j �MQ�M��l���E�    �E������E�   ��Uă��UċM諛���E������E� �E�    �E�    �	�Eȃ��EȋM�;M�(  �	�UЃ��UЋEЋM�A��t�EЋM�A�   k� �E�;�t�ʋU�R�M��a��� ��t�M�Q�M���`���UЉU��   �E�EĉEЋMЋU�J�   k� �M�;�t�EЋM�A��u.�}�s�EĉE���E�   �M�Q�M��`���U���EȉE��\�MQ�UR�#`��������u�MЋU�4J�M蠅����;�t(�}�s�MĉM���E�   �U�R�M��>`���M����E�������Uυ�t�EP�MQ�_�����Ѕ�t��q����E��E��E������M��Lf���E��M�d�    Y^�M�3���v����]����������������������������������������������������������������������������������������������������������������������������������������������������������U����M��E��H(��t�U�B�E��	�M�Q�U��E���,Pj �M�Q�V�����U��B�E�H.��v	�E��a�	�U�B �E�M���,Qj �U�R��U�����M��A�U�B/��v	�E��	�M�Q$�U��E���,Pj �M�Q�U�����U��B�E���,Pj �   k� �E�H�R��q�����M�f�A�U���,Rj �   k� �U�B�Q�q�����U�f�B��]� �������������������������������������������������������������������������������U��Q�M��EPj �   k� �E��R�#q�����M�f�A�URj �   k� �U�B�Q��p�����U�f�B��]�4 ������������������������������������U���4���3ŉE�VW�M̍E�P�M蘈���}̃��   ���M̃�Qj �M�V��P�)T�����ỦB�Ẽ�Pj �M�$S��P�	T�����M̉A�Ũ�Rj hX���S�����M̉A_^�M�3���s����]� ��������������������������������������������������U����M��E��H(��t�U�B8�E��	�M�Q<�U��E�P�O�����M��A�U�B.��v	�E�p��	�M�QH�U�E�P�uO�����M��A�U�B/��v	�E�t��	�M�QL�U��E�P�EO�����M��A�   k� �M�Q@�M�f�f�Q�   k� �U�BD�U�f�f�B��]� ��������������������������������������������������������������U��Q�M��   k� �U�B0�U�f�f�B�   k� �E�H4�E�f�
f�H��]�4 �����������������U���4���3ŉE�VW�M̍E�P�M�h����}̃��   ���M��~��P�8N�����M̉A�M�_��P�!N�����ỦBhЦ�N�����M̉A_^�M�3���q����]� ���������������������������������������������U��Q3��E��E���]�����������������U��Q3��E��E���]�����������������U��Q�E�M���E��]��������������U��Q�E�M���E��]��������������U��Q�E�M���E��]��������������U��Q�E�M���E��]��������������U��Q�E�M���E��]��������������U��Q�E���]������U��Q�E���]������U��E]���������U��E]���������U�����E���E�M���M�U;Ut8�E;Et0�M��E�;�}����M��U��M�;�}�   �4뮋E;Et	�E�������M;Mt	�E�   ��E�    �U��U��E���]�������������������������������������������������U��EP�MQ�UR�EP�MQ������]����������������U��Q�E+E���E��M+M��9M�w!�U���R�EP�M+M����Q�UR�\�����E���]�����������������������������U��EP�MQ�UR�EP�MQ�-�����]����������������U���3�f�E��E�    �MQ�U�Rj�EP�M�Q�������f�E���]����������������������������U���3�f�E��E�    �MQ�U�Rj�EP�M�Q讝����f�E���]����������������������������U���,�E�    �EP�y�������E�M�M��E�    �U�U���E�+E�E��M�M�M�U����U��}� v)�EP�M�Q�U�R�E�P�M�Q�������E�}� �붋U����U�h  hЕ�>���P3ɋE��   �������Q��L�����E؋E؉E��M��M��E�    �$�U�+U�U��EE�E�M����M��U���U�}� v)�EP�M�Q�U�R�EP�M�Q�z������E�}� ��3ҋE�f��E���]������������������������������������������������������������������������������������U���,�E�    �EP� x�������E�M�M��E�    �U�U���E�+E�E��M�M�M�U����U��}� v)�EP�M�Q�U�R�E�P�M�Q蚛�����E�}� �붋U����U�h�  hЕ辁��P3ɋE��   �������Q�lK�����E؋E؉E��M��M��E�    �$�U�+U�U��EE�E�M����M��U���U�}� v)�EP�M�Q�U�R�EP�M�Q��������E�}� ��3ҋE�f��E���]������������������������������������������������������������������������������������U��Q�E���]������U��Q�E���]������U��E]���������U��E]���������U��E]���������U��j�hx�d�    P��`���3�P�E�d�    �M��E�   ���̉eȍEP�!]���E�M�M��E����̉e��UR�]���E�E�E��E��M�Q�M��N���E�U�U��E����̉e��E�P聘���E܋M܉M��E��U�R�M��c\���E؋E؉E��E����̉e��U�R�J����E��E��M��C����EЋEЉE��E��M��P���E��M��P���E� �M�P���E������M��O���E̋M�d�    Y��]� �������������������������������������������������������������������������������������U��j�h��d�    P��`���3�P�E�d�    �M��E�   ���̉eȍEP��}���E�M�M��E����̉e��UR�}���E�E�E��E��M�Q�M���V���E�U�U��E����̉e��E�P�P���E܋M܉M��E��U�R�M��m����E؋E؉E��E����̉e��U�R��O���E��E��M��c���EЋEЉE��E��M��	W���E��M���V���E� �M��V���E������M��V���E̋M�d�    Y��]� �������������������������������������������������������������������������������������U��Q�M��EP�b�����P�MQ�U�R�\�������]� ����������������������U��j�h1�d�    P�����3�P�E�d�    �M�EPj�g�����E��E�    �}� t�MQ�������U�� ��M��M���E�    �U�U��E������M�d�    Y��]� ������������������������������������������U��EP�v�����P�MQ�M�~��]�������������������U��Q�M��EP譌����P�MQ�U�R�jU������]� ����������������������U��j�hq�d�    P�����3�P�E�d�    �M�EPj�f�����E��E�    �}� t�MQ�.������U�� ��M��M���E�    �U�U��E������M�d�    Y��]� ������������������������������������������U��EP�������P�MQ�M�E\��]�������������������U��Q�E;Eu�M�U��E�A�E�{�yhQ  h ��MQ�UR�a����hR  h ��EP�R�����MQ�UR�pA�����E��E�P�MQ�UR�EP�n����P�MQ�n����P�UR��{�����E��]���������������������������������������������������U��Q�E;Eu�M�U��E�A�E�{�yhQ  h ��MQ�UR��`����hR  h ��EP�]������MQ�UR�	d�����E��E�P�MQ�UR�EP��m����P�MQ�m����P�UR�b�����E��]���������������������������������������������������U��Q�M��EP�M�Q�/D������]� �������������������U��Q�M���]� ���U��EP�M��V��]����������������U��Q�M��EP�M�Q�<|������]� �������������������U��Q�M���]� ���U��EP�M�'L��]����������������U��E]���������U��E]���������U��E]���������U��E]���������U��j�h��d�    P��$���3�P�E�d�    j �M��P���E�    �H��E���L���E�M�Q�M��s���E�}� t�n�}� t�U��U��`�EP�M�Q��b�������uhDq�M��U��hPP�U�R��v���.�E��E�M��H��U��U�E��M�B�ЋM�Q�d������U�U��E������M��{���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��IO���E�    ���E���aK���E�M�Q�M�r���E�}� t�n�}� t�U��U��`�EP�M�Q�d�������uhDq�M��^T��hPP�U�R�u���.�E��E�M����U��U�E��M�B�ЋM�Q�$������U�U��E������M���y���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M��	N���E�    �(��E����!J���E�M�Q�M�Yq���E�}� t�n�}� t�U��U��`�EP�M�Q�Uc�������uhDq�M��S��hPP�U�R�Dt���.�E��E�M��(��U��U�E��M�B�ЋM�Q��~�����U�U��E������M��x���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h8�d�    P��$���3�P�E�d�    j �M���L���E�    ����E����H���E�M�Q�M�p���E�}� t�n�}� t�U��U��`�EP�M�Q�hZ�������uhDq�M���Q��hPP�U�R�s���.�E��E�M�����U��U�E��M�B�ЋM�Q�}�����U�U��E������M��Vw���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hh�d�    P��$���3�P�E�d�    j �M��K���E�    ����E����G���E�M�Q�M��n���E�}� t�n�}� t�U��U��`�EP�M�Q��O�������uhDq�M��P��hPP�U�R��q���.�E��E�M�����U��U�E��M�B�ЋM�Q�d|�����U�U��E������M��v���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��IJ���E�    ����E���aF���E�M�Q�M�m���E�}� t�n�}� t�U��U��`�EP�M�Q�Y�������uhDq�M��^O��hPP�U�R�p���.�E��E�M�����U��U�E��M�B�ЋM�Q�${�����U�U��E������M���t���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��	I���E�    �,��E����!E���E�M�Q�M�Yl���E�}� t�n�}� t�U��U��`�EP�M�Q�fz�������uhDq�M��N��hPP�U�R�Do���.�E��E�M��,��U��U�E��M�B�ЋM�Q��y�����U�U��E������M��s���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M���G���E�    ����E����C���E�M�Q�M�k���E�}� t�n�}� t�U��U��`�EP�M�Q�/\�������uhDq�M���L��hPP�U�R�n���.�E��E�M�����U��U�E��M�B�ЋM�Q�x�����U�U��E������M��Vr���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h(�d�    P��$���3�P�E�d�    j �M��F���E�    �0��E����B���E�M�Q�M��i���E�}� t�n�}� t�U��U��`�EP�M�Q�h�������uhDq�M��K��hPP�U�R��l���.�E��E�M��0��U��U�E��M�B�ЋM�Q�dw�����U�U��E������M��q���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hX�d�    P��$���3�P�E�d�    j �M��IE���E�    � ��E���aA���E�M�Q�M�h���E�}� t�n�}� t�U��U��`�EP�M�Q�l3�������uhDq�M��^J��hPP�U�R�k���.�E��E�M�� ��U��U�E��M�B�ЋM�Q�$v�����U�U��E������M���o���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��	D���E�    �4��E����!@���E�M�Q�M�Yg���E�}� t�n�}� t�U��U��`�EP�M�Q�
^�������uhDq�M��I��hPP�U�R�Dj���.�E��E�M��4��U��U�E��M�B�ЋM�Q��t�����U�U��E������M��n���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M���B���E�    ���E����>���E�M�Q�M�f���E�}� t�n�}� t�U��U��`�EP�M�Q�2�������uhDq�M���G��hPP�U�R�i���.�E��E�M����U��U�E��M�B�ЋM�Q�s�����U�U��E������M��Vm���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��A���E�    �<��E����=���E�M�Q�M��d���E�}� t�n�}� t�U��U��`�EP�M�Q豄�������uhDq�M��F��hPP�U�R��g���.�E��E�M��<��U��U�E��M�B�ЋM�Q�dr�����U�U��E������M��l���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M��I@���E�    �8��E����a<���E�M�Q�M�c���E�}� t�n�}� t�U��U��`�EP�M�Q��l�������uhDq�M��^E��hPP�U�R�f���.�E��E�M��8��U��U�E��M�B�ЋM�Q�$q�����U�U��E������M���j���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hH�d�    P��$���3�P�E�d�    j �M��	?���E�    ���E���!;���E�M�Q�M�Yb���E�}� t�n�}� t�U��U��`�EP�M�Q�O�������uhDq�M��D��hPP�U�R�De���.�E��E�M����U��U�E��M�B�ЋM�Q��o�����U�U��E������M��i���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hx�d�    P��$���3�P�E�d�    j �M���=���E�    ���E����9���E�M�Q�M�a���E�}� t�n�}� t�U��U��`�EP�M�Q��F�������uhDq�M���B��hPP�U�R�d���.�E��E�M����U��U�E��M�B�ЋM�Q�n�����U�U��E������M��Vh���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��<���E�    ���E���8���E�M�Q�M��_���E�}� t�n�}� t�U��U��`�EP�M�Q�^�������uhDq�M��A��hPP�U�R��b���.�E��E�M����U��U�E��M�B�ЋM�Q�dm�����U�U��E������M��g���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��I;���E�    ����E���a7���E�M�Q�M�^���E�}� t�n�}� t�U��U��`�EP�M�Q�Ql�������uhDq�M��^@��hPP�U�R�a���.�E��E�M�����U��U�E��M�B�ЋM�Q�$l�����U�U��E������M���e���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M��	:���E�    � ��E����!6���E�M�Q�M�Y]���E�}� t�n�}� t�U��U��`�EP�M�Q�4�������uhDq�M��?��hPP�U�R�D`���.�E��E�M�� ��U��U�E��M�B�ЋM�Q��j�����U�U��E������M��d���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h8�d�    P��$���3�P�E�d�    j �M���8���E�    ����E����4���E�M�Q�M�\���E�}� t�n�}� t�U��U��`�EP�M�Q�+�������uhDq�M���=��hPP�U�R�_���.�E��E�M�����U��U�E��M�B�ЋM�Q�i�����U�U��E������M��Vc���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hh�d�    P��$���3�P�E�d�    j �M��7���E�    �$��E����3���E�M�Q�M��Z���E�}� t�n�}� t�U��U��`�EP�M�Q�!B�������uhDq�M��<��hPP�U�R��]���.�E��E�M��$��U��U�E��M�B�ЋM�Q�dh�����U�U��E������M��b���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��I6���E�    ����E���a2���E�M�Q�M�Y���E�}� t�n�}� t�U��U��`�EP�M�Q�H�������uhDq�M��^;��hPP�U�R�\���.�E��E�M�����U��U�E��M�B�ЋM�Q�$g�����U�U��E������M���`���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��	5���E�    �@��E����!1���E�M�Q�M�YX���E�}� t�n�}� t�U��U��`�EP�M�Q�6(�������uhDq�M��:��hPP�U�R�D[���.�E��E�M��@��U��U�E��M�B�ЋM�Q��e�����U�U��E������M��_���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M���3���E�    ���E����/���E�M�Q�M�W���E�}� t�n�}� t�U��U��`�EP�M�Q��J�������uhDq�M���8��hPP�U�R�Z���.�E��E�M����U��U�E��M�B�ЋM�Q�d�����U�U��E������M��V^���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h(�d�    P��$���3�P�E�d�    j �M��2���E�    �D��E����.���E�M�Q�M��U���E�}� t�n�}� t�U��U��`�EP�M�Q�,�������uhDq�M��7��hPP�U�R��X���.�E��E�M��D��U��U�E��M�B�ЋM�Q�dc�����U�U��E������M��]���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hX�d�    P��$���3�P�E�d�    j �M��I1���E�    ���E���a-���E�M�Q�M�T���E�}� t�n�}� t�U��U��`�EP�M�Q�K^�������uhDq�M��^6��hPP�U�R�W���.�E��E�M����U��U�E��M�B�ЋM�Q�$b�����U�U��E������M���[���E܋M�d�    Y��]��������������������������������������������������������������������������U��Q�M��EP�M���L���E���]� ��������������������U��Q�M��M��a���E���]�����������U��Q�M��EP�M��L���E���]� ��������������������U��Q�M��M��@a���E���]�����������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��F���E�    �M��t��U��E�B(�MQ�UR�M��f7���E������E��M�d�    Y��]� �����������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��xE���E�    �M��L��U��E�B(�MQ�UR�M��+���E������E��M�d�    Y��]� �����������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��M��F���E�    �M���d���E������E��M�d�    Y��]� ������������������������U��j�h�d�    PQ���3�P�E�d�    �M��M��g���E�    �M���e���E������E��M�d�    Y��]� ������������������������U��Q�M��EP�M���G���M��U�B�A�E���]� ������������������������U��j�hH�d�    PQ���3�P�E�d�    �M��M��Fn���E�    �EP�M���Y���M��U�Q�E������E��M�d�    Y��]� ���������������������������U��Q�M��M���m���E��@    �E���]�����������������U��Q�M��EP�M��+���M��U�B�A�E���]� ������������������������U��j�hx�d�    PQ���3�P�E�d�    �M��M��l\���E�    �EP�M���X���M��U�Q�E������E��M�d�    Y��]� ���������������������������U��Q�M��M��\���E��@    �E���]�����������������U��Q�M��EP�M��l���E���]� ��������������������U��Q�M��EP�MQ�M���)���E���]� ����������������U��Q�M��EP�M��$���E���]� ��������������������U��Q�M��EP�MQ�M��j���E���]� ����������������U��Q�M��M��S���E��@    �M��A    �E���]�����������������������U��Q�M��M���R���E��@    �M��A    �E���]�����������������������U��Q�M��EP�M��Tk���E���]� ��������������������U��Q�M��M��mI���E���]�����������U��Q�M��EP�M���U���E���]� ��������������������U��Q�M��M��qO���E���]�����������U��Q�M��E���]� ����������������U��Q�M��E���]�������������������U��Q�M��E���]� ����������������U��Q�M��E���]�������������������U����M��E�P�M���P�M�����j j �M��_���MQ�^����P�M��S���E���]� ������������������������U��j�h��d�    P�����3�P�E�d�    �M�E�P�M�Q�M������^��P�M��a���E�    j j �M��t^���P�Rj �EP�M��[���E������E�M�d�    Y��]� �������������������������������������U��j�h��d�    P�����3�P�E�d�    �M�M��LG��P�M������E�    j j �M���]���EP�MQ�M��"���E������E�M�d�    Y��]� ����������������������������������������U��j�h�d�    P�����3�P�E�d�    �M�M��F��P�M�� ���E�    j j �M��3]���EP�M��;g���E������E�M�d�    Y��]� �����������������������������U��j�h8�d�    P�����3�P�E�d�    �M�M��F��P�M�����E�    j j �M��\���EP�MQ�M���"���E������E�M�d�    Y��]� �����������������������������������������U��j�hh�d�    P�����3�P�E�d�    �M�M��|E��P�M������E�    j j �M��\���E������E�M�d�    Y��]����������������������������U����M��E�P�M��!��P�M�����j j �M���7���MQ�����P�M��h3���E���]� ������������������������U��j�h��d�    P�����3�P�E�d�    �M�E�P�M�Q�M�N!�����
^��P�M��G���E�    j j �M��Q7�����Rj �EP�M��'$���E������E�M�d�    Y��]� �������������������������������������U��j�h��d�    P�����3�P�E�d�    �M�M��@J��P�M�����E�    j j �M��6���EP�MQ�M��y/���E������E�M�d�    Y��]� ����������������������������������������U��j�h��d�    P�����3�P�E�d�    �M�M��I��P�M�����E�    j j �M��6���EP�M��^���E������E�M�d�    Y��]� �����������������������������U��j�h(�d�    P�����3�P�E�d�    �M�M��I��P�M��v���E�    j j �M��5���EP�MQ�M��TL���E������E�M�d�    Y��]� �����������������������������������������U��j�hX�d�    P�����3�P�E�d�    �M�M��pH��P�M������E�    j j �M���4���E������E�M�d�    Y��]����������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��R*���E�    �M��ĝ�UR�M��VK���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M���)���E�    �M�����UR�M���a���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M���0���E�    �M����UR�M��_���E������E��M�d�    Y��]� ���������������������������������������U��j�h�d�    PQ���3�P�E�d�    �M��EP�M��E0���E�    �M��̟�UR�M���U���E������E��M�d�    Y��]� ���������������������������������������U��j�hH�d�    PQ���3�P�E�d�    �M��EP�M���<���E�    �M��D��UR�M��0���E������E��M�d�    Y��]� ���������������������������������������U��j�hx�d�    PQ���3�P�E�d�    �M��EP�M��1<���E�    �M�����UR�M��*O���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��W���E�    �M����UR�M�� ���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M���V���E�    �M����UR�M��_+���E������E��M�d�    Y��]� ���������������������������������������U��j�h�d�    PQ���3�P�E�d�    �M��EP�M��u-���E�    �M��8��UR�M������E������E��M�d�    Y��]� ���������������������������������������U��j�h8�d�    PQ���3�P�E�d�    �M��EP�M���,���E�    �M����UR�M������E������E��M�d�    Y��]� ���������������������������������������U��j�hh�d�    PQ���3�P�E�d�    �M��EP�M��U,���E�    �M��X��UR�M�����E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M���+���E�    �M��0��UR�M������E������E��M�d�    Y��]� ���������������������������������������U��Q�M��EPj�MQ�UR�M���&���E�� ���E���]� ����������������U��Q�M��EPj �MQ�UR�M��&���E�� ���E���]� ����������������U��Q�M��EPj�MQ�UR�M��5���E�� ̠�E���]� ����������������U��Q�M��EPj �MQ�UR�M��y5���E�� ���E���]� ����������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��5*���E�    �M��@��UR�M��;X���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��)���E�    �M����UR�M��61���E������E��M�d�    Y��]� ���������������������������������������U��j�h(�d�    PQ���3�P�E�d�    �M��EP�M��)���E�    �M�����UR�M��0���E������E��M�d�    Y��]� ���������������������������������������U��j�hX�d�    PQ���3�P�E�d�    �M��EP�M��(���E�    �M��d��UR�M��]H���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M���'���E�    �M��ġ�UR�EP�M���+���E������E��M�d�    Y��]� ����������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��e'���E�    �M�����UR�EP�M��3���E������E��M�d�    Y��]� ����������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M�����E�    �M��4��UR�M��@J���E������E��M�d�    Y��]� ���������������������������������������U��j�h�d�    PQ���3�P�E�d�    �M��EP�M������E�    �M����UR�M��T���E������E��M�d�    Y��]� ���������������������������������������U��j�hS�d�    PQ���3�P�E�d�    �M��EP�M��%���E�    �M��h�j �M����4���E��UR�M��M$���E������E��M�d�    Y��]� ��������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��%���E�    �M��Оj �M����4���E��UR�M��	���E������E��M�d�    Y��]� ��������������������������������������U��Q�M��E��M��E���]� ��������U��Q�M��EP�M��t$���M�����E���]� �����������U��Q�M��EP�M��D$���M�����E���]� �����������U��Q�M��EP�M��$���M�����E���]� �����������U��Q�M��M��g"����]��������������U��Q�M��M��G"����]��������������U��Q�M��E�� t��M��l3���M��A����]�������������U��Q�M��E�� L��M������M������]�������������U��Q�M��M��GG���M�� ����]����������������������U��Q�M��M��l$���M������]����������������������U��Q�M��M���J����]��������������U��Q�M��M��x6����]��������������U��Q�M��M������]��������������U��Q�M��M��	����]��������������U��Q�M��M������]��������������U��Q�M��M�������]��������������U��Q�M�j j�M��lH���M�������]������������������U��Q�M�j j�M��y$���M��i����]������������������U��Q�M��E�� ĝ�M���&����]���������������������U��Q�M��E�� ���M���&����]���������������������U��Q�M��E�� ��M��QR�J�����M�������]����������������������U��Q�M��E�� ̟�M��QR�LJ�����M������]����������������������U��Q�M��E�� D��M��y t�U��BP�J�����M��QR��I�����M������]������������������������������U��Q�M��E�� ���M��y t�U��BP�I�����M��QR�I�����M��6����]������������������������������U��Q�M��E�� ��M��,1����]���������������������U��Q�M��E�� ��M���0����]���������������������U��Q�M��E�� 8��M��U����]���������������������U��Q�M��E�� ��M��%����]���������������������U��Q�M��E�� X��M�������]���������������������U��Q�M��E�� 0��M�������]���������������������U��Q�M��E�� ���M��i<����]���������������������U��Q�M��E�� ���M��9<����]���������������������U��Q�M��E�� ̠�M��	����]���������������������U��Q�M��E�� ���M��	����]���������������������U��Q�M��E�� @��M�������]���������������������U��Q�M��E�� ��M������]���������������������U��Q�M��E�� ���M��u����]���������������������U��Q�M��E�� d��M��E����]���������������������U��Q�M��E�� ġ�M��M"���M������]�������������U��Q�M��E�� ���M��>���M�������]�������������U��Q�M��E�� 4��M��@���M��E����]�������������U��Q�M��E�� ��M������M��dE����]�������������U��Q�M��E�� h��M����H���M��J����]����������U��Q�M��E�� О�M�����G���M������]����������U��Q�M��E��Q�E������]��������U��Q�M��M�������]��������������U��Q�M��M������]��������������U��Q�M��E�� ���M������]���������������������U��Q�M��EP�M�����E���]� ��������������������U��Q�M��EP�M�����E���]� ��������������������U��Q�M��EP�M��Q/���M��U�B�A�E���]� ������������������������U��Q�M��EP�M��p���M��U�B�A�E���]� ������������������������U����M��E��;Mtv�M�� ���} th�U�U��E����t�U����U���E����E��M�+M�M�h-  h�j�U�R�������M���U��: t�E�P�MQ�U��P�������E���]� ����������������������������������������������U����M��E�;E��   j j�M��n@��3�t�U�R�M�Z���P�M���*���E�P�M�E���P�M�Q�M��8���P�<5�����Ѕ�t,���ĉe�P�M� �����̉e�Q�M����M���?����UR�?����P�M��4���E���]� ���������������������������������������������������U����M��E�;EtZ�M�Q�M����P�U�R�M�����P�4��������t%3�t!j j�M��e?���U�R�M�U���P�M���)���EP�M�� ���E���]� ��������������������������������������������U����M��E�;E��   j j�M��+��3�t�U�R�M����P�M�����E�P�M����P�M�Q�M�����P��)�����Ѕ�t,���ĉe�P�M�������̉e�Q�M�<���M��)����UR������P�M��C���E���]� ���������������������������������������������������U����M��E�;EtZ�M�Q�M�)��P�U�R�M����P�)��������t%3�t!j j�M��"���U�R�M����P�M�����EP�M��� ���E���]� ��������������������������������������������U����M��E��x t4�MQ�U��J���f�E��[-��f�E��E�P�M�Q�������Ѕ�t�E�� �E���]� ���������������������������U����M��E��x t4�MQ�U��J�� ��f�E���B��f�E��E�P�M�Q�y=�����Ѕ�t�E�� �E���]� ���������������������������U��Q�M��E��M���E�     �E���]� �������������U����M��EP�M��G2���M��U�A;Bu	�E�   ��E�    �E���]� ��������������������U����M��EP�M��H"���M��U�A;Bu	�E�   ��E�    �E���]� ��������������������U����M��EP�M��-���ȅ�u	�E�   ��E�    �E���]� ���������������������������U����M��EP�M���C���ȅ�u	�E�   ��E�    �E���]� ���������������������������U��Q�M��E��H;Msh�  h �h,��
�����M������U�P��]� �������������������U��Q�M��E��H;Msh�  h �h,��^
�����M��W���U�P��]� �������������������U��Q�M��E��H;Msh�  h �h,��
�����M���'���U�P��]� �������������������U��Q�M��E��H;Msh�  h �h,��	�����M��6'���U�P��]� �������������������U��QV�M��M�������tG�E��x t>�M�������
���M�9Ar'�M�������
�����M�����P�V�M�;Aw_jOh �h�o�(	������i��t3�u#hjhpjj jPh �j��������u�j jPh �h`�h�k��5�����U��B^��]������������������������������������������������������������U��QV�M��M�������tG�E��x t>�M�������O&���M�9Ar'�M�������8&�����M�����P�V�M�;Aw_jOh �h�o�(������i��t3�u#hjhpjj jPh �j��������u�j jPh �h�h�k��4�����U��B^��]������������������������������������������������������������U��Q�M��M������]��������������U��Q�M��M��3����]��������������U��Q�M��E��H��u�M��k����U��: uh�  h��h �������E�f�@��]�����������������������������U��Q�M��E��H��u�M���7���U��: uh�  h��h �������E�f�@��]�����������������������������U��Q�M��E���]�������������������U��Q�M��E���]�������������������U��QV�M��M�������t0�E��x t'�M��r������c�����M��a����H�N�E�;Pw_jmh �h���������i��t3�u#hjhpjj jnh �j���������u�j jnh �hh�h�k�2�����M��Q���E��P�E�^��]�������������������������������������������������������U��QV�M��M�������t0�E��x t'�M��������#�����M��q����H�N�E�;Pw_jmh �h��������i��t3�u#hjhpjj jnh �j��������u�j jnh �hh�h�k�1�����M��Q���E��P�E�^��]�������������������������������������������������������U��Q�M��E��8 uh  h��hh��Q�����M���'���E���]����������������������������U��Q�M��E��8 uh  h��hh�������M������E���]����������������������������U��Q�M��E���]� ����������������U��Q�M��E���]�������������������U��Q�M��E���]� ����������������U��Q�M��E���]�������������������U��Q�M��EP�M��)���M��U�A+B����]� ���������U��Q�M��EP�M�����M��U�A+B����]� ���������U��j�h��d�    P�����3�P�E�d�    �M��E�    �E�P�M������E�    �MQ�M����P�M�����U����U��E������M��o����E�M�d�    Y��]� ���������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M��EP�M�Q�M���<���E�U�U��E�    �M���3���E��E������M������E�M�d�    Y��]� ������������������������������������������U��j�h(�d�    P�����3�P�E�d�    �M��E�    �E�P�M���"���E�    �MQ�M��S���P�M��"���U����U��E������M������E�M�d�    Y��]� ���������������������������������������������U��j�hX�d�    P�����3�P�E�d�    �M��EP�M�Q�M������E�U�U��E�    �M��"-���E��E������M��6����E�M�d�    Y��]� ������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M��E�    �E�P�M��V����E�    �MQ�M�����P�M�:����U����U��E������M�������E�M�d�    Y��]� ���������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M��E�    �E�P�M��� ���E�    �MQ�M��!��P�M�� ���U����U��E������M������E�M�d�    Y��]� ���������������������������������������������U��QV�M��M��'�����tW�E��x tN�M��Q�E�4B�M������������;�r/�M����������������M�������H�N�E��H�E�A;�shh�   h �h��u�������i��t3�u&hjhpjj h�   h �j�d�������u�j h�   h �h��h�k�+�����U��B�M�H�E��P�E�^��]� �����������������������������������������������������������������U��QV�M��M��������tW�E��x tN�M��Q�E�4B�M���������s��;�r/�M���������`�����M������H�N�E��H�E�A;�shh�   h �h��E�������i��t3�u&hjhpjj h�   h �j�4�������u�j h�   h �hp�h�k��)�����U��B�M�H�E��P�E�^��]� �����������������������������������������������������������������U��Q�M��EP�M�������E���]� ��������������������U��Q�M��EP�M���3���E���]� ��������������������U��Q�M��EP�M��������]� �������U��Q�M��EPj�M��5����]� ��������������������U��Q�M��EP�M��.�����]� �������U��Q�M��EPj�M��:����]� ��������������������U��Q�M��E��P�M��9 ����]� ���������������������U��Q�M��E��P�M������]� ���������������������U��Q�M��M��"���E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q�O������E���]� ��������������������U��Q�M��M������E��t�M�Q�������E���]� ��������������������U��Q�M��M��x����E��t�M�Q��������E���]� ��������������������U��Q�M��M������E��t�M�Q�������E���]� ��������������������U��Q�M��M�����E��t�M�Q�O������E���]� ��������������������U��Q�M��M��|����E��t�M�Q�������E���]� ��������������������U��Q�M��M�������E��t�M�Q��������E���]� ��������������������U��Q�M��M��Z ���E��t�M�Q�������E���]� ��������������������U��Q�M��M��
����E��t�M�Q�O������E���]� ��������������������U��Q�M��M������E��t�M�Q�������E���]� ��������������������U��Q�M��M���4���E��t�M�Q��������E���]� ��������������������U��Q�M��M��@���E��t�M�Q�������E���]� ��������������������U��Q�M��M��^���E��t�M�Q�O������E���]� ��������������������U��Q�M��M��4����E��t�M�Q�������E���]� ��������������������U��Q�M��M��/ ���E��t�M�Q��������E���]� ��������������������U��Q�M��M��5���E��t�M�Q�������E���]� ��������������������U��Q�M��M�����E��t�M�Q�O������E���]� ��������������������U��Q�M��M�����E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q��������E���]� ��������������������U��Q�M��M��-���E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q�O������E���]� ��������������������U��Q�M��M��{����E��t�M�Q�������E���]� ��������������������U��Q�M��M��>���E��t�M�Q��������E���]� ��������������������U��Q�M��M��.���E��t�M�Q�������E���]� ��������������������U��Q�M��M��v����E��t�M�Q�O������E���]� ��������������������U��Q�M��M��! ���E��t�M�Q�������E���]� ��������������������U��Q�M��M��&���E��t�M�Q��������E���]� ��������������������U��Q�M��M��U���E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q�O������E���]� ��������������������U��Q�M��M��E&���E��t�M�Q�������E���]� ��������������������U����M��M������j�M������M���M����P�U��P�M������M���E����]����������������������������U����M��M�����j�M��y���M���M����P�U��P�M�����M���E����]����������������������������U����M��E�xs"�M�Q��R�E��P�M���Q������+�U��R�E���P�M�Q�M���������<���U�B    �E��M�Q�P�E��M�Q�Pj j �M�"����]� ���������������������������������������U����M��E�xs"�M�Q��R�E��P�M���Q��������+�U��R�E���P�M�Q�M��8������K���U�B    �E��M�Q�P�E��M�Q�Pj j �M�)�����]� ���������������������������������������U����M��E��8 t
�M���U��	�E����E��E���]����������������������U��Q�M���]� ���U��Q�M���]� ���U��Q�M��}u�EP�M������M�HR�������� �EP�MQ�M�������U�PP��������]� ��������������������������������U��Q�M��}u�EP�M��R���M�HR�&����� �EP�MQ�M��0���U�PP��������]� ��������������������������������U��QV�M��M��G�����t�M��;������M�1���;�thh�   h �hh����������m��t3�u&h(nhpjj h�   h �j���������u�j h�   h �h��h�o�v����^��]� ���������������������������������������U��QV�M��M�������t�M��{������M�q���;�thh�   h �hh���������m��t3�u&h(nhpjj h�   h �j��������u�j h�   h �h��h�o�����^��]� ���������������������������������������U��j�h��d�    PQ�� SVW���3�P�E�d�    �e��M�E���E�M����;E�s�M�M��R�E�3ҹ   ��U�J��;�w�8�U�r��M�����+ƋM�9Aw�U�B��M�A�E���M�����E��E�    �U�R�M��I����E܋E��P�M��$����E؋M؉M��g�e��U�U��E��E�P�M������EԋM��Q�M�������EЋUЉU��j j�M�����j j ����J��E�   ��E�   �/J��E�������E������} v�EP�M��w���P�M�Q������j j�M�����U�R�E��P�M�Q�M��s����������U�E�B�MQ�M������M�d�    Y_^[��]� ������������������������������������������������������������������������������������������������������������������������U��j�h�d�    PQ�� SVW���3�P�E�d�    �e��M�E���E�M������;E�s�M�M��R�E�3ҹ   ��U�J��;�w�8�U�r��M�����+ƋM�9Aw�U�B��M�A�E���M��{����E��E�    �U�R�M��4����E܋E��P�M������E؋M؉M��g�e��U�U��E��E�P�M�������EԋM��Q�M��]����EЋUЉU��j j�M������j j �j���IL��E�   ��E�   �_L��E�������E������} v�EP�M�����P�M�Q�Q�����j j�M������U�R�E��P�M�Q�M��^������q���U�E�B�MQ�M������M�d�    Y_^[��]� ������������������������������������������������������������������������������������������������������������������������U������3ŉE��M��E�    �E��P�M�Q�UR�E�P�=&������t�M�M���   k� �L�M�E�M�3�������]� ���������������������������U������3ŉE��M��E�    �E��P�M�Q�UR�E�P�%������t�M�M���   k� �L�M�E�M�3��>�����]� ���������������������������U����M��E�    �E��P�M�Qj�UR�E�P�%������}���  f�M��f�U�f�U�f�E���]� ����������������������������������U����M��E�    �E��P�M�Qj�UR�E�P�$������}���  f�M��f�U�f�U�f�E���]� ����������������������������������U����M��E��8 u	�E�   ��E�    �E���]�������������������������U����M�3�f�E��M��U�Q�E�P�M��+����M�HR��������]� �����������������������U����M�3�f�E��M��U�Q�E�P�M�����M�HR�[�������]� �����������������������U����E�E�M��%�U���U�E�� t�M��+�U���U�E��t�M��#�U���U�E�� .�M���M�U��*�E���E��M��t�U�E��M���M�U�� 0  �U��E��tP�}�    u�E�f�.�}� 0  u�E�A��}�   u�E�E��E�G�M��M��U��U��E�M���U���U��N�}�    u�E�f�.�}� 0  u�E�a��}�   u�E�e��E�g�E��E��M��M��U�E���M���M�U�� �E��]����������������������������������������������������������������������������������U����E�E�M��%�U���U�E�� t�M��+�U���U�E��t�M��#�U���U�E�� .�M���M�U��*�E���E��M��t�U�E��M���M�U�� 0  �U��E��tP�}�    u�E�f�.�}� 0  u�E�A��}�   u�E�E��E�G�M��M��U��U��E�M���U���U��N�}�    u�E�f�.�}� 0  u�E�a��}�   u�E�e��E�g�E��E��M��M��U�E���M���M�U�� �E��]����������������������������������������������������������������������������������U��j�hf�d�    P���   ���3ŉE�VP�E�d�    h`  hx��EP�4������}0 v�M ���+t�E ���-u	�E�   ��E�    �U��U��M�	��% 0  = 0  tǅ|��� ��Jǅ|���$��E���;E0w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M���|���R�   k� M Q�Z�����E�f�(�f�U��i����   k� � �   k� ��T��   k� �T�R�   k� M Q������E���`���R�M������l�����l�����\����E�    ��\���Q� �����E��E�������`����M���j0�M��g���f�E�j �U0R�M��6����E�   j �M��,���P�E E0P�   k� U R�M��D����p���P�M������d�����d�����h����E���h���R�P������E��E���p��������E�P�M��u����E��M�����f�E��M$�M��U�;U0u �E�E��E��M�Q�U$R�E�P�M������e�M�M��M��U�R�E,P�M�Q�M�����U�R�E(P�M���Q�M�����M����f���U�R�M��3���f�0�E�P�M$Q�U�R�M��e��j �M������E��E����tY�U����~O�M���E�+E�;�s?�M���E�+E��M�Qj�U�R�M�����   �� �M����~	�E����E�뜍M������E0�M�l�����t�����x�����x��� |(	��t��� v�M�D���;E0v�M�7���+E0�E���E�    �M��M��M����%�  �E��}�@ty�}�   tp�U�R�EP�MQ�UR��<���P�MQ��������@�U�E�E�    �M�Qj �M������P�UR�EP��T���Q�UR�[�������P�M�U�   �}�   um�E�Pj �M�����P�MQ�UR��,���P�MQ��������@�U�E�M�Q�UR�EP�MQ��D���R�EP�!������P�M�U�E�    �5�E�Pj �M��:���P�MQ�UR��4���P�MQ��������@�U�E�M0+M�Q�U�R�M�� ���P�EP�MQ��L���R�EP�q�������P�M�Uj j �M�����E�P�MQ�UR�EP�MQ�UR�q�����E��M��(����E������M��1����E�M�d�    Y^�M�3��������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P���   ���3ŉE�VP�E�d�    h`  hx��EP�������}0 v�M ���+t�E ���-u	�E�   ��E�    �U��U��M�)��% 0  = 0  tǅ|��� ��Jǅ|���$��E���;E0w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M���|���R�   k� M Q�z�����E�f�(�f�U������   k� � �   k� ��T��   k� �T�R�   k� M Q�-�����E���`���R�M�������l�����l�����\����E�    ��\���Q�������E��E�������`����m���j0�M����f�E�j �U0R�M��/���E�   j �M�����P�E E0P�   k� U R�M��B�����p���P�M�4�����d�����d�����h����E���h���R�z������E��E���p���������E�P�M�������E��M������f�E��M$�M��U�;U0u �E�E��E��M�Q�U$R�E�P�M�������e�M�M��M��U�R�E,P�M�Q�M�������U�R�E(P�M���Q�M�������M������f���U�R�M������f�0�E�P�M$Q�U�R�M�����j �M�������E��E����tY�U����~O�M���E�+E�;�s?�M���E�+E��M�Qj�U�R�M��@����   �� �M����~	�E����E�뜍M��E���E0�M������t�����x�����x��� |(	��t��� v�M�d���;E0v�M�W���+E0�E���E�    �M��M��M����%�  �E��}�@ty�}�   tp�U�R�EP�MQ�UR��<���P�MQ�E������@�U�E�E�    �M�Qj �M��|���P�UR�EP��T���Q�UR��������P�M�U�   �}�   um�E�Pj �M��9���P�MQ�UR��,���P�MQ�X�������@�U�E�M�Q�UR�EP�MQ��D���R�EP�������P�M�U�E�    �5�E�Pj �M������P�MQ�UR��4���P�MQ���������@�U�E�M0+M�Q�U�R�M�����P�EP�MQ��L���R�EP��������P�M�Uj j �M�����E�P�MQ�UR�EP�MQ�UR�������E��M��H����E������M�������E�M�d�    Y^�M�3��������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��M������M��%����E��Q�M��~���j�U��P�M�����M��    ��]�����������������������������U����M��M������M�������E��Q�M�����j�U��P�M��K���M��    ��]�����������������������������U��Q�M��M�.����E��]� ��������U��Q�M��M�t����E��]� ��������U��j�hT�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h^  hЕ�M�Qj4�-������E��E�    �}� t:j �M����P�M��9����E��U��U��E��E����E��M�Q�M�����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��e���   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �m����E�hs  hЕ�M�Qj4��������E��E�    �}� t:j �M�Y���P�M�������E��U��U��E��E����E��M�Q�M��.���E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��%���   �M�d�    Y��]��������������������������������������������������������������������������U��j�hM�d�    P��x���3ŉE�P�E�d�    �E�    �} ��   �E�8 ��   �*����E�jCh ��M�Qj�������E��E�    �}� tbj �U�R�M������E��E��E��E��MЃ��MЋM�����P��|��������E��U��U��E�   �EЃ��EЋM�Q�M������E���E�    �UȉU��E�   �E�M���E�   �UЃ�t�e����|����	���E������EЃ�t�e���M������   �M�d�    Y�M�3�������]������������������������������������������������������������������������������������������U��j�h��d�    P��x���3ŉE�P�E�d�    �E�    �} ��   �E�8 ��   �����E�jCh ��M�Qj�������E��E�    �}� tbj �U�R�M�R����E��E��E��E��MЃ��MЋM������P��|���������E��U��U��E�   �EЃ��EЋM�Q�M��I	���E���E�    �UȉU��E�   �E�M���E�   �UЃ�t�e����|�������E������EЃ�t�e���M��m����   �M�d�    Y�M�3�������]������������������������������������������������������������������������������������������U��j�hT�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�hO  hЕ�M�QjD�m������E��E�    �}� t:j �M�����P�M��y����E��U��U��E��E����E��M�Q�M��N����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�hl
  hЕ�M�QjD�-������E��E�    �}� t:j �M����P�M��9����E��U��U��E��E����E��M�Q�M��9����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��e���   �M�d�    Y��]��������������������������������������������������������������������������U��j�h1�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �m����E�jMh���M�Qj��������E��E�    �}� t:j �M�\���P�M�������E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��(���   �M�d�    Y��]�����������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �-����E�jMh���M�Qj�������E��E�    �}� t:j �M����P�M������E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]�����������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�h�  h��M�Qj�m������E��E�    �}� t:j �M�����P�M��y����E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]��������������������������������������������������������������������������U��j�hd�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h�  h��M�Qj�-������E��E�    �}� t:j �M����P�M��9����E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��e ���   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �m����E�h�  h��M�Qj��������E��E�    �}� t:j �M�Y���P�M�������E��U��U��E��E����E��M�Q�M��Ͷ���E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��%����   �M�d�    Y��]��������������������������������������������������������������������������U��j�hD�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �-����E�h�  h��M�Qj�������E��E�    �}� t:j �M����P�M������E��U��U��E��E����E��M�Q�M�蠻���E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�h(  h��M�QjX�m������E��E�    �}� t<jj �M�����P�M��w����E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]������������������������������������������������������������������������U��j�h$�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h(  h��M�QjX�-������E��E�    �}� t<jj �M����P�M��7����E��U��U��E��E����E��M�Q�M��8����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��c����   �M�d�    Y��]������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �m����E�h(  h��M�QjX��������E��E�    �}� t<jj �M�W���P�M�������E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��#����   �M�d�    Y��]������������������������������������������������������������������������U��j�h�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �-����E�h(  h��M�QjX譿�����E��E�    �}� t<jj �M����P�M������E��U��U��E��E����E��M�Q�M��7����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�������   �M�d�    Y��]������������������������������������������������������������������������U��j�ht�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�h  h`��M�Qj�m������E��E�    �}� t:j �M�����P�M��y����E��U��U��E��E����E��M�Q�M��2����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h  h`��M�Qj�-������E��E�    �}� t:j �M����P�M��9����E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��e����   �M�d�    Y��]��������������������������������������������������������������������������U��j�hT�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �m����E�hD  h`��M�Qj�������E��E�    �}� t:j �M�Y���P�M�������E��U��U��E��E����E��M�Q�M��W����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��%����   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �-����E�hD  h`��M�Qj譺�����E��E�    �}� t:j �M����P�M������E��U��U��E��E����E��M�Q�M��y����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h4�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�h�   h`��M�Qj�m������E��E�    �}� t<jj �M�����P�M��w����E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h�   h`��M�Qj�-������E��E�    �}� t<jj �M����P�M��7����E��U��U��E��E����E��M�Q�M�藽���E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��c����   �M�d�    Y��]������������������������������������������������������������������������U��j�h�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �m����E�h�   h|��M�QjD�������E��E�    �}� t:j �M�Y���P�M�������E��U��U��E��E����E��M�Q�M��T����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��%����   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �-����E�h�   h|��M�QjD譵�����E��E�    �}� t:j �M����P�M������E��U��U��E��E����E��M�Q�M�褭���E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�h  h|��M�Qj�m������E��E�    �}� t:j �M�����P�M��y����E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�hd�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h|  h|��M�Qj�-������E��E�    �}� t:j �M����P�M��9����E��U��U��E��E����E��M�Q�M��0����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��e����   �M�d�    Y��]��������������������������������������������������������������������������U����M������E�U��E�M��U��P�E��]� ���������������������U��Q�M�������]�����������������U����M������E��}� t�E�P�M����o����M�Q�������M����1����Ѕ�u�M����ҳ���E���E�h��E��]�������������������������������U��j�h��d�    P��   ���3ŉE�VP�E�d�    �M�q���% 0  = 0  u%�EP�MQ�UR�EP�MQ�UR���������  ��L���P�M������\�����\�����T����E�    ��T���R���������p����E�������L����N����E�P��p��������E�   �M�M��E� ��P���R�M�>�����X�����X�����`����E���`���Q�)�������h����E���P��������U�R�   k�����Q�   k� ��P��h���������MQ�UR�p���������t�h�M�����Ⱥ   k��T�;�u�E�� +�M����M��M�k����3�M�ݸ���и   k�
�D�;�u�M��-�U����U��M�6����E� �E�    �E�    j �M�躨����|�����|������t��|��������   ��E��M������MQ�UR����������te�M�D�����Q�U�R�'������E��}�
sD�}�$|�E����E��.�}� u�}� u� �M��U�������M����M��U����U��x����;  �M��װ����u3�f��v������p�������f��v���f��v���f��x���j j�M��U����E��E�    ��M�����UR�EP�������ȅ���   �M�g�����R�E�P�J������E��}�
s~�E��}�$|�M����M��.�}� u�}� u� �U��E������
�U����U��E����E��M�Q�M���������t%�E�P�M�謥����l�����l��������l�����M�M�Q�M�腥�����t!��x�����t�M誶������x���;�t��j j�M�訳���E����E�������}� u�"�M�Q�M��+������~�E����E���E��M�����   �}� ��   ��|������u�{�t�M����M�t��|����2�E�P�M��ͤ���;�u"�}� u"��|����2�E�P�M�諤���;�}�E��%�   �� ��|������~��|�������|����_����E��M�������E���t�}� u�M��0�U����U��EP�MQ�������Ѕ�tE�M�k�������p����P�����;�u(�j����   k� � �M����E����E��M�����}� uj��E��M�����MQ�UR�<���������t'�M������Ⱥ   k� �T�;�u�E����E�붃}� }�M��0�U����U��E����E���E��M�4����MQ�UR�����������tI�M葴����Q�U�R�t������E��}�
s(�}�$} �E��M�������E����E��M����M���U�����  �EP�MQ�f������Ѕ���  �M�!������   k��L�;�t �M�����и   k��D�;��i  �M��e�U����U��M�Z����E� �E�    �EP�MQ�������Ѕ�t�h�M誳�����   k��L�;�u�U��+�E����E��M�����3�M�u����Ⱥ   k�
�T�;�u�E�� -�M����M��M������UR�EP�l������ȅ�t*�M�+����и   k� �D�;�u�E��M������M���t�U��0�E����E���E��M�h����MQ�UR����������tI�M�Ų����Q�U�R�������E��}�
s(�}�} �E��M�������E����E��M����M���U���u�E���u�M�M��U�� �E���d����E������M��j�����d����M�d�    Y^�M�3�������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h6�d�    P��   ���3ŉE�VP�E�d�    �M����% 0  = 0  u%�EP�MQ�UR�EP�MQ�UR蕬������  ��L���P�M�M�����\�����\�����T����E�    ��T���R萓������p����E�������L��������E�P��p����Ү���E�   �M�M��E� ��P���R�M�޹����X�����X�����`����E���`���Q�1�������h����E���P���腒���U�R�   k���إQ�   k� إP��h����w����MQ�UR�(���������t�h�M�����Ⱥ   k��T�;�u�E�� +�M����M��M�m����3�M�x����и   k�
�D�;�u�M��-�U����U��M�8����E� �E�    �E�    j �M��Z�����|�����|������t��|��������   ��E��M������MQ�UR����������te�M�������Q�U�R��������E��}�
sD�}�$|�E����E��.�}� u�}� u� �M��U���إ��M����M��U����U��x����;  �M��w�����u3�f��v������p�������f��v���f��v���f��x���j j�M�������E��E�    ��M�����UR�EP�������ȅ���   �M������R�E�P��������E��}�
s~�E��}�$|�M����M��.�}� u�}� u� �U��E���إ�
�U����U��E����E��M�Q�M��`������t%�E�P�M��L�����l�����l��������l�����M�M�Q�M��%������t!��x�����t�M�E�������x���;�t��j j�M��H����E����E�������}� u�"�M�Q�M��˚�����~�E����E���E��M�����   �}� ��   ��|������u�{�t�M����M�t��|����2�E�P�M��m����;�u"�}� u"��|����2�E�P�M��K����;�}�E��%�   �� ��|������~��|�������|����_����E��M��a����E���t�}� u�M��0�U����U��EP�MQ�������Ѕ�tE�M��������p����&�����;�u(�
����   k� � �M����E����E��M�����}� uj��E��M�����MQ�UR蝫��������t'�M薾���Ⱥ   k� �T�;�u�E����E�붃}� }�M��0�U����U��E����E���E��M�6����MQ�UR�3���������tI�M�,�����Q�U�R�(������E��}�
s(�}�$} �E��M���إ��E����E��M����M���U�����  �EP�MQ�Ǫ�����Ѕ���  �M輽�����   k��L�;�t �M蠽���и   k��D�;��i  �M��e�U����U��M�\����E� �E�    �EP�MQ��������Ѕ�t�h�M�E������   k��L�;�u�U��+�E����E��M�����3�M�����Ⱥ   k�
�T�;�u�E�� -�M����M��M������UR�EP�ͩ�����ȅ�t*�M�Ƽ���и   k� �D�;�u�E��M������M���t�U��0�E����E���E��M�j����MQ�UR�g���������tI�M�`�����Q�U�R�\������E��}�
s(�}�} �E��M���إ��E����E��M����M���U���u�E���u�M�M��U�� �E���d����E������M��
�����d����M�d�    Y^�M�3�赭����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P���   ���3ŉE�VP�E�d�    ��0���P�M�&�����@�����@�����8����E�    ��8���R�_�������T����E�������0����ǈ���E�P��T����{����E�   ��4���Q�M�������<�����<�����D����E���D���P謻������L����E���4����h����M�Q�   k��P�   k� ���R��L����|����E��x���ƅw��� �MQ�UR����������t�z�M腤���Ⱥ   k��T�;�u"��x���� +��x�������x����M�ն���<�M�G����и   k��D�;�u ��x����-��x�������x����M藶����x���� 0��x�������x�����x����x��x�������x���ƅ��� ǅp���    ǅd���    �MQ�UR����������u�M詣���Ⱥ   k� �T�;�t�e�EP�M����P�������ȅ�tB�M�o����и   k��D�;�t�M�S����Ⱥ   k��T�;�u
�M軵���ƅ���j �M��H�����`�����`������t��`��������   �ƅ����M�r����MQ�UR������������   �M�ˢ����Q�U�R��������h�����h���se��p���$|��d�������d����F��h��� u��p��� u�2��x�����h���������x�������x�����p�������p����J����  �M��7�����u3�f��Z������T�������f��Z���f��Z���f��\���j j�M�赛���E�ǅl���    ��M�k����UR�EP�	������ȅ��.  �M�ġ����R�E�P��������h�����h�����   ƅ�����p���$|��d�������d����F��h��� u��p��� u�2��x�����h�������
��x�������x�����p�������p�����l���Q�M��������t(��l���P�M��Տ����P�����P��������P�����V��l���Q�M�諏�����t!��\�����t�M�Р������\���;�t�"�j j�M��Ν����l�������l���������l��� u�.��l���Q�M��E������~��l�������l����ƅw�����w�������   ��l��� ��   ��`������u
�   �   ��l�������l���t��`����2��l���P�M��Ɏ���;�u(��l��� u(��`����2��l���P�M�衎���;�}	ƅw����%�   �� ��`������~��`�������`����A����E��M�贔���������t!��p��� u��x����0��x�������x����EP�MQ�������Ѕ�tN�M�O�������T����4�����;�u1�N����   k� � ��x�������x�������x����M荱����p��� ��   �ƅ����M�o����MQ�UR����������t-�M�̞���Ⱥ   k� �T�;�u��d�������d���뭃�d��� }'��x����0��x�������x�����d�������d����ƅ����M�����MQ�UR����������tg�M�G�����Q�U�R�*�������h�����h���s@��p���$}2��x�����h���������x�������x�����p�������p����s�����������  �EP�MQ��������Ѕ���  �M趝�����   k��L�;�t �M蚝���и   k��D�;���  ��x����p��x�������x����M����ƅ��� ǅp���    �EP�MQ莨�����Ѕ�t�z�M�0������   k��L�;�u"��x����+��x�������x����M耯���<�M�����Ⱥ   k��T�;�u ��x���� -��x�������x����M�B����UR�EP��������ȅ�t-�M蟜���и   k� �D�;�uƅ����M� �����������t��x����0��x�������x����ƅ����M�ʮ���MQ�UR�h���������tg�M�'�����Q�U�R�
�������h�����h���s@��p���}2��x�����h���������x�������x�����p�������p����s�����w�����u�������u	�M��x�����x���� �E��d����ǅH���    �E������M�薐����H����M�d�    Y^�M�3��A�����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P���   ���3ŉE�VP�E�d�    ��0���P�M�&�����@�����@�����8����E�    ��8���R�i|������T����E�������0�����{���E�P��T���諗���E�   ��4���Q�M�������<�����<�����D����E���D���P�~������L����E���4����h{���M�Q�   k���P�   k� �¤�R��L����Z����E��x���ƅw��� �MQ�UR�����������t�z�M耫���Ⱥ   k��T�;�u"��x���� +��x�������x����M�7����<�M�B����и   k��D�;�u ��x����-��x�������x����M�������x���� 0��x�������x�����x����x��x�������x���ƅ��� ǅp���    ǅd���    �MQ�UR����������u�M褪���Ⱥ   k� �T�;�t�e�EP�M�m���P�q������ȅ�tB�M�j����и   k��D�;�t�M�N����Ⱥ   k��T�;�u
�M�����ƅ���j �M��H�����`�����`������t��`��������   �ƅ����M�Ծ���MQ�UR�і����������   �M�Ʃ����Q�U�R�´������h�����h���se��p���$|��d�������d����F��h��� u��p��� u�2��x�����h����������x�������x�����p�������p����J����  �M��7�����u3�f��Z������T�����|��f��Z���f��Z���f��\���j j�M�赎���E�ǅl���    ��M�ͽ���UR�EP�ʕ�����ȅ��.  �M迨����R�E�P軳������h�����h�����   ƅ�����p���$|��d�������d����F��h��� u��p��� u�2��x�����h��������
��x�������x�����p�������p�����l���Q�M��������t(��l���P�M��Ղ����P�����P��������P�����V��l���Q�M�諂�����t!��\�����t�M�˧������\���;�t�"�j j�M��ΐ����l�������l���������l��� u�.��l���Q�M��E������~��l�������l����ƅw�����w�������   ��l��� ��   ��`������u
�   �   ��l�������l���t��`����2��l���P�M��Ɂ���;�u(��l��� u(��`����2��l���P�M�衁���;�}	ƅw����%�   �� ��`������~��`�������`����A����E��M�贇���������t!��p��� u��x����0��x�������x����EP�MQ�Q������Ѕ�tN�M�J�������T����j�����;�u1�N����   k� � ��x�������x�������x����M������p��� ��   �ƅ����M�Ѻ���MQ�UR�Β��������t-�M�ǥ���Ⱥ   k� �T�;�u��d�������d���뭃�d��� }'��x����0��x�������x�����d�������d����ƅ����M�L����MQ�UR�I���������tg�M�B�����Q�U�R�>�������h�����h���s@��p���$}2��x�����h����������x�������x�����p�������p����s�����������  �EP�MQ輑�����Ѕ���  �M豤�����   k��L�;�t �M蕤���и   k��D�;���  ��x����p��x�������x����M�H���ƅ��� ǅp���    �EP�MQ�~�����Ѕ�t�z�M�+������   k��L�;�u"��x����+��x�������x����M�����<�M�����Ⱥ   k��T�;�u ��x���� -��x�������x����M褸���UR�EP衐�����ȅ�t-�M蚣���и   k� �D�;�uƅ����M�b�����������t��x����0��x�������x����ƅ����M�,����MQ�UR�)���������tg�M�"�����Q�U�R��������h�����h���s@��p���}2��x�����h����������x�������x�����p�������p����s�����w�����u�������u	�M��x�����x���� �E��d����ǅH���    �E������M�薃����H����M�d�    Y^�M�3��A�����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hh�d�    P�����3�P�E�d�    �M��E�P�M�-����E�M�M��E�    �U�R�!������E��E������M���n���	�E(���E(�M(�����   �E(���%uO�U(���U(j �E(�Q�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M���M��B$�Ћ�P�M�U�   �E(��� uB��M�V����UR�EP��������ȅ�t�M賊����RjH�M��(�������t���<j �M萊����Q�M��'����ЋE(�;�t�U ����M ����M���������UR�EP薕�����ȅ�t�U ����M ��U�E��M�J�E�M�d�    Y��]�$ �����������������������������������������������������������������������������������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M��E�P�M�����E�M�M��E�    �U�R�io�����E��E������M���l���	�E(���E(�M(�����   �E(���%uO�U(���U(j �E(�Q�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M���M��B$�Ћ�P�M�U�   �E(��� uB��M蘱���UR�EP蕉�����ȅ�t�M莜����RjH�M�軉������t���<j �M�k�����Q�M��]q���ЋE(�;�t�U ����M ����M�$��������UR�EP�v�����ȅ�t�U ����M ��U�E��M�J�E�M�d�    Y��]�$ �����������������������������������������������������������������������������������������������������������������������U��j�h��d�    P���   ���3ŉE�VP�E�d�    �EP�J�������X����M�Q��X����x����E�    �M�������u3�f��f������X����ʤ��f��f���f��f���f��h����MQ蚝������8����U�R�   k���`�Q�   k� `�P��8����y����M��|����UR�EP�������ȅ�t�z�M艆���и   k��D�;�u"��|����+��|�������|����M�٘���<�M�K������   k��L�;�u ��|����-��|�������|����M蛘���M��   �M�}   uǅ`���   �I�}   uǅD���   �(�} uǅL���    �
ǅL���
   ��L�����D�����D�����`�����`�����p����E� ƅw��� �UR�EP踵�����ȅ���   �M�s����и   k� �D�;���   �E��M�ӗ���MQ�UR�q���������tb�M�0����Ⱥ   k��T�;�t�M�������   k��L�;�u*��p��� t	��p���uǅp���   �E� �M�\������p��� u
ǅp���   ��p��� t6��p���
t-��p���uǅT���   �
ǅT���   ��T�����H����
ǅH���
   ��H�����@����M�Qj�M��~���E�ǅx���    �   k�E��<�����M躖���MQ�UR�X����������!  �M������Q�U�R���������P�����P���;�@�����   ��|�����P�����`����w�����u��|������0t$��|���;�<���s��|�������|���ƅw����E���x���P�M��Hr�����t(��x���R�M��1r����\�����\��������\����
�V��x���P�M��r�����t!��h�����t�M�,�������h���;�t�"�j j�M��*�����x�������x���������x��� u�+��x���P�M��q�����~��x�������x�����E� j �M���r����l����E�����   ��x��� ��   ��l������u
�   �   ��x�������x���t��l����1��x���R�M��q��� ;�u(��x��� u%��l����1��x���R�M���p��� ;�}�E� �%�   �� ��l����
��~��l�������l����G����U���t%��w�����u��|����0��|�������|�����E���u	�M��|�����|���� ��p�����4����E� �M��v���E������M��v����4����M�d�    Y^�M�3��R�����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h �d�    P���   ���3ŉE�VP�E�d�    �EP�c������X����M�Q��X�������E�    �M��}x����u3�f��f������X����g��f��f���f��f���f��h����MQ�be������8����U�R�   k�����Q�   k� ��P��8����v���M��|����UR�EP�_m�����ȅ�t�z�M�����и   k��D�;�u"��|����+��|�������|����M蛧���<�M覒�����   k��L�;�u ��|����-��|�������|����M�]����M��   �M�}   uǅ`���   �I�}   uǅD���   �(�} uǅL���    �
ǅL���
   ��L�����D�����D�����`�����`�����p����E� ƅw��� �UR�EP��~�����ȅ���   �M�Α���и   k� �D�;���   �E��M蕦���MQ�UR�~��������tb�M苑���Ⱥ   k��T�;�t�M�o������   k��L�;�u*��p��� t	��p���uǅp���   �E� �M�������p��� u
ǅp���   ��p��� t6��p���
t-��p���uǅT���   �
ǅT���   ��T�����H����
ǅH���
   ��H�����@����M�Qj�M��uv���E�ǅx���    �   k�E��<�����M�|����MQ�UR�y}���������!  �M�n�����Q�U�R�j�������P�����P���;�@�����   ��|�����P����������w�����u��|������0t$��|���;�<���s��|�������|���ƅw����E���x���P�M��j�����t(��x���R�M��j����\�����\��������\����
�V��x���P�M��gj�����t!��h�����t�M臏������h���;�t�"�j j�M��x����x�������x���������x��� u�+��x���P�M��j�����~��x�������x�����E� j �M��>k����l����E�����   ��x��� ��   ��l������u
�   �   ��x�������x���t��l����1��x���R�M��{i��� ;�u(��x��� u%��l����1��x���R�M��Si��� ;�}�E� �%�   �� ��l����
��~��l�������l����G����U���t%��w�����u��|����0��|�������|�����E���u	�M��|�����|���� ��p�����4����E� �M��o���E������M��o����4����M�d�    Y^�M�3������]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���@���3ŉE��E܉EԋMQ�UR�c���������t�[j �M�x����Q�M �z���E��Uۃ�+u�E�� +�Mԃ��MԋM�X���� �Uۃ�-u�E�� -�Mԃ��MԋM�6����E� �UR�EP�Ч�����ȅ�t,j �M�w����R�M �$z������0u�E��M������Mڅ�t�U��0�Eԃ��EԹ   k��D܉E���E��M軉���MQ�UR�Y���������tFj �M�w����Q�M �y���E��Uۃ�0|$�Eۃ�9�MԊUۈ�E�;E�s	�Mԃ��M���Uڅ�u�E܉EԋM�� �E�    �U�Rj
�E�P�M�Q�4������E��E�    �UR�EP�܁�����ȅ�t	�UЃ��UЍE�9E�t�}� u�M�;M|�U;U�}�EЃ��E���M�Ủ�EЋM�3��"|����]����������������������������������������������������������������������������������������������������������������������������������U���@���3ŉE��E܉EԋMQ�UR��c��������t�[j �M�~�����Q�M �p^���E��Uۃ�+u�E�� +�Mԃ��MԋM�:���� �Uۃ�-u�E�� -�Mԃ��MԋM�����E� �UR�EP�v�����ȅ�t,j �M������R�M ��]������0u�E��M�ӝ����Mڅ�t�U��0�Eԃ��EԹ   k��D܉E���E��M蝝���MQ�UR�u��������tFj �M葈����Q�M �]���E��Uۃ�0|$�Eۃ�9�MԊUۈ�E�;E�s	�Mԃ��M���Uڅ�u�E܉EԋM�� �E�    �U�Rj
�E�P�M�Q�}�����E��E�    �UR�EP�tb�����ȅ�t	�UЃ��UЍE�9E�t�}� u�M�;M|�U;U�}�EЃ��E���M�Ủ�EЋM�3��y����]����������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P���  ���3ŉE�VP�E�d�    ��t���ǅ|���    h�  h��E�HQ�R�E�HQ�R��������E��tQ������Q�M�h}���������������� ����E�    �� ���P�x������p����E������������	V���O������Q�M�}���������������������E�   ������P�ܜ������p����E������������U��ƅ���� ƅw��� �M������E�   ��4���Q��p����a���M�������E�������R�M�|���������������������E�������Q�x�������$����E��������4U���UR�   k�����Q�   k� ��P��$����H���ǅ`���    ���`�������`������������K  ��`����>  ��`�����4�����<�����<����� ��<�����<���X�	  ��<��������$����U�R��p��������E�������R���E��M������u=�EP�MQ��������Ѕ�t&�M�p�����M��{��� ;�tj �M��v���Q��`���uH�M��X�����w;�MQ�UR��{��������u�M�fp�����M��2{���;�t
j �M���u����h���R�M�� h���������������������E�������Q������p���E���h�����[���������/����M�s����UR�EP�������ȅ�tv��\���R�M��Y��������������x����E���|�������|�����x���R�������������t)�M�o����������h���;�uǅ(���   �
ǅ(���    ��(�����^����E�   ��|�����t��|������\����
[����^�����t������D���R�M��WX���������������������E�	������Q������5�����\����E���D����Z����\�����tƅ�����E��������Z���E��M���d���  �EP�MQ��y�����Ѕ�t�t  ������P��p����Q���������������������E�
��|�������|����������
�����vej ������P��p�����P���������������������E�   ��|�������|����������h���0�M��m����;�uǅ���   �
ǅ���    �������Z����E�
   ��|�����t��|������������c���E�   ��|�����t��|�����������c����Z�����t?�M����������R��p�����O��������������P�M��e���������bc���!  �����Q��p����|���������������������E���|�������|���������跞����vej ������Q��p����q|���������������������E�   ��|�������|����������0g���0�M�l����;�uǅ���   �
ǅ���    �������S����E�   ��|�����t��|��������xb���E�   ��|�����t��|����������Tb����S�����tF�M�~����H���P��p����{��������������Q�M��Ed����H����b��ƅw�����   ��,���R��p����_N���������������|�����uǅ ���   �
ǅ ���    �� �����_�����,����a����_�����t�f������R��p�����z��������������������uǅ,���   �
ǅ,���    ��,�����[����������Na����[�����tƅw�����  ǅT���    ��p�����k����8�����d���R��p����%����E���d�����c����u3�f��B������p�����t��f��B���f��B���f��H�����H�����t��d����Y��� ��|e��M��|���MQ�UR蔚��������t?�M�Sj����Q�UR�6�������h�����h���
s��h�������Q�M��aY����M  j j�M���c���E�ǅx���    ��M�w|���UR�EP�������ȅ���   �M��i����R�EP賜������h�����h���
sW��h�������R�M���X����x���P�M��MX�����t(��x���R�M��6X���������������������
�K��x���P�M��X�����t�M�<i������H���;�t�"�j j�M��:f����x�������x���������x��� u�.��x���R�M��W��� ��~��x�������x����ƅ������d�����W����L�������������   ��x��� ��   ��L������u
�   �   ��x�������x���t��L����0��x���Q�M��$W���;�u(��x��� u(��L����0��x���Q�M���V���;�}	ƅ�����%�   �� ��L������~��L�������L����A�����������t �E��M��]���E���d�����\����  �E��M���\����p����ɞ��f��D����UR�EP�ڗ�����ȅ���   ��D�������   �M�g������D���;���   �UR�M��y��P著��������t\��T���;�8���}N�M�Bg����R�EP�%�������h�����h���
s'��h�������R�M��PV����T�������T���눋�T���;�8���}ƅ�����M���_����u	ƅ�����+���T�������T�����T���;�8���}j0�M���U�����E���d����[���   ��`���u�vƅo��� ��M��x���MQ�UR虖��������t)�M�Xf����QjH��$����ʒ���Ѕ�t	ƅo���븋�`�����4����� u��o�����uƅ������������������  �M��ė������  �������G���E���,���Q�M��]���������������������E�������P�������f���E���,����zQ����M�x����P���Q�M���N����������������|����E���|����� ��|�����|���Q������耂�����z���Ѕ�t@�EP�MQ�\������Ѕ�t)�M�e�����������^��� ;�uǅ0���   �
ǅ0���    ��0�����]����E�   ��|����� t��|���ߍ�P����P����]�����t������8���Q�M���M���������������������E�������P��������y����g����E���8����FP����g�����tƅ�����E��������pP����������tj �M��̉�����w�����tj-jj �M��d����M�Q�M�X����|�����@��|����E��M��Y���E������M��Z���E�M�d�    Y^�M�3��i����]� ����������z�  �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P���  ���3ŉE�VP�E�d�    ��t���ǅ|���    h�  h��E�HQ�R�E�HQ�R�X{�����E��tQ������Q�M�xi���������������� ����E�    �� ���P�4�������p����E������������B���O������Q�M�'i���������������������E�   ������P�7M������p����E�������������A��ƅ���� ƅw��� �M��s���E�   ��4���Q��p����H����M������E�������R�M�h���������������������E�������Q��C������$����E��������DA���UR�   k���P�Q�   k� P�P��$����6U��ǅ`���    ���`�������`������������K  ��`����>  ��`�����4�����<�����<����� ��<�����<���X�	  ��<��������$����U�R��p�����^���E�������^���E��M������u=�EP�MQ��]�����Ѕ�t&�M��p�����M���w��� ;�tj �M��
����Q��`���uH�M�诈����w;�MQ�UR��J��������u�M�qp�����M��w���;�t
j �M�跆����h���R�M�躃���������������������E�������Q�������V���E���h����aP���������t����M�����UR�EP��\�����ȅ�tv��\���R�M��O��������������x����E���|�������|�����x���R������g_������t)�M�o��������������;�uǅ(���   �
ǅ(���    ��(�����^����E�   ��|�����t��|������\����O����^�����t������D���R�M���N���������������������E�	������Q������^����\����E���D����)O����\�����tƅ�����E�������W<���E��M��Qm���  �EP�MQ��H�����Ѕ�t�t  ������P��p����l���������������������E�
��|�������|����������a�����vej ������P��p����Jl���������������������E�   ��|�������|����������j���0�M��m����;�uǅ���   �
ǅ���    �������Z����E�
   ��|�����t��|�����������Kl���E�   ��|�����t��|�����������'l����Z�����t?�M�X���������R��p����vk��������������P�M��-O����������k���!  �����Q��p����_���������������������E���|�������|���������������vej ������Q��p����g_���������������������E�   ��|�������|����������h���0�M�l����;�uǅ���   �
ǅ���    �������S����E�   ��|�����t��|���������j���E�   ��|�����t��|�����������j����S�����tF�M������H���P��p����^��������������Q�M���M����H����j��ƅw�����   ��,���R��p�����i���������������Ӄ����uǅ ���   �
ǅ ���    �� �����_�����,����/j����_�����t�f������R��p�����]���������������r�����uǅ,���   �
ǅ,���    ��,�����[�����������i����[�����tƅw�����  ǅT���    ��p���������8�����d���R��p�����R���E���d�����O����u3�f��B������p���訁��f��B���f��B���f��H�����H�����t��d����E��� ��|e��M�h���MQ�UR�eW��������t?�M�^j����Q�UR�Zu������h�����h���
s��h�����P�Q�M��qE����M  j j�M���O���E�ǅx���    ��M��~���UR�EP��V�����ȅ���   �M��i����R�EP��t������h�����h���
sW��h�����P�R�M���D����x���P�M��]D�����t(��x���R�M��FD���������������������
�K��x���P�M��D�����t�M�Gi������H���;�t�"�j j�M��JR����x�������x���������x��� u�.��x���R�M���C��� ��~��x�������x����ƅ������d�����C����L�������������   ��x��� ��   ��L������u
�   �   ��x�������x���t��L����0��x���Q�M��4C���;�u(��x��� u(��L����0��x���Q�M��C���;�}	ƅ�����%�   �� ��L������~��L�������L����A�����������t �E��M��I���E���d����I����  �E��M���H����p����c��f��D����UR�EP�T�����ȅ���   ��D�������   �M�g������D���;���   �UR�M�^|��P�bT��������t\��T���;�8���}N�M�Mg����R�EP�Ir������h�����h���
s'��h�����P�R�M��`B����T�������T���눋�T���;�8���}ƅ�����M���K����u	ƅ�����+���T�������T�����T���;�8���}j0�M���A�����E���d�����G���   ��`���u�vƅo��� ��M�m{���MQ�UR�jS��������t)�M�cf����QjH��$����S���Ѕ�t	ƅo���븋�`�����4����� u��o�����uƅ������������������  �M��~������  �������
S���E���,���Q�M��Ny���������������������E�������P�������gL���E���,�����E����M�z����P���Q�M��PE����������������|����E���|����� ��|�����|���Q��������u�����U���Ѕ�t@�EP�MQ�-R�����Ѕ�t)�M�&e�����������u��� ;�uǅ0���   �
ǅ0���    ��0�����]����E�   ��|����� t��|���ߍ�P����E����]�����t������8���Q�M��rD���������������������E�������P�������NT����g����E���8�����D����g�����tƅ�����E���������1����������tj �M���u�����w�����tj-jj �M��t����M�Q�M��D����|�����@��|����E��M��E���E������M��b���E�M�d�    Y^�M�3��U����]� ����u���w�j�  �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��4���E��}� t�E�P�M�����>���M�Q�yw�����M����j���Ѕ�u�M����2D���E���E�К�E��]�������������������������������U��Q�M��E�� ��]�����������������U����M��E��H�9 t�U��B,��M���E�    �E����]�����������������U����M��E��H�9 t�U��B,��M���E�    �E����]�����������������U����M��E��H,����E��H,��U��B��M��U��B����U��B��E���]��������������������������������U����M��E��H,����E��H,��U��B��M��U��B����U��B��E���]��������������������������������U����M��M��X��;Es�M��gm���E��H;Ms�U��BP�MQ�M��s4���J�U��t2�}s,�E��M;Hs�U�U��	�E��H�M��U�Rj�M��ir����} u
j �M���V���} v	�E�   ��E�    �E��]� �����������������������������������������U����M��M��F*��;Es�M���|���E��H;Ms�U��BP�MQ�M��ZO���J�U��t2�}s,�E��M;Hs�U�U��	�E��H�M��U�Rj�M���M����} u
j �M���@���} v	�E�   ��E�    �E��]� �����������������������������������������U����E�ŝ��E� �E�ŝ��E�    �	�E����E��M�;Ms�UU��3E��E�iM�� �M��ԋE���]��������������������������U����E�E��M��%�U����U��E�� t�M��+�U����U��E��t�M��#�U����U��   k� �U�
��Lt�   k� �E��M���E����E��-�M��I�U����U��E�� 6�M����M��U��4�E����E��M��   �M�}�   u�E�o�:�}�   t�   �� �E��M���U��t�E�X��E�x�E��E��M��M��U��E���M����M��U�� �E��]��������������������������������������������������������������������������������������U����E�E��M��%�U����U��E�� t�M��+�U����U��E��t�M��#�U����U��   k� �U�
��Lt�   k� �E��M���E����E��-�M��I�U����U��E�� 6�M����M��U��4�E����E��M��   �M�}�   u�E�o�:�}�   t�   �� �E��M���U��t�E�X��E�x�E��E��M��M��U��E���M����M��U�� �E��]��������������������������������������������������������������������������������������U����M��E��8 t.�M��	�v��f�E���]��f�E��U�R�E�P�(�����ȅ�t�U��    �E��@��M��A ��]�������������������������������������U����M��E��8 t.�M��	�h��f�E��6s��f�E��U�R�E�P��m�����ȅ�t�U��    �E��@��M��A ��]�������������������������������������U��j�h@�d�    PQ��@���3ŉE�SVWP�E�d�    �e��M��E�P�M�k]���}���,�   ���M�M_���E��M��A    �U��B    �E��@    �M��A    �E�    �U���,Rj �E��HQ��6�����E��U��E��B�M�Qj �M��Q=����M��U��j j ��\�������E�������E������U��B(��t�M��Q(�U��	�E��H)�M��U��E��P�M��y |	�U��z|
�E��@    �M��Q.R�E��H*Q�U��B+P�M��� Q�M��-0���U��B/P�M��Q,R�E��H-Q�U���$R�M��0���E��t,jhȦ�M��� Q�\2����jhȦ�U���$R�F2�����M�d�    Y_^[�M�3��G����]� �������������������������������������������������������������������������������������������������������������������������U��j�hp�d�    PQ��@���3ŉE�SVWP�E�d�    �e��M��E�P�M�+[���}���,�   ���M�]���E��M��A    �U��B    �E��@    �M��A    �E�    �U���,Rj �E��HQ�4�����E��U��E��B�M�Qj �M��a@����M��&:��j j �Z������E�������E������U��B(��t�M��Q(�U��	�E��H)�M��U��E��P�M��y |	�U��z|
�E��@    �M��Q.R�E��H*Q�U��B+P�M��� Q�M��Qo���U��B/P�M��Q,R�E��H-Q�U���$R�M��*o���E��t,jhȦ�M��� Q�0����jhȦ�U���$R�0�����M�d�    Y_^[�M�3��lE����]� �������������������������������������������������������������������������������������������������������������������������U���4���3ŉE�VW�M̍E�P�M�Y���}̃��   ���_^�M�3��D����]� ������������������������������U���4���3ŉE�VW�M̍E�P�M�X���}̃��   ���_^�M�3��QD����]� ������������������������������U����M��E�P�M��i����P�E��H�P��]� �����������������������U����M��E�P�M�i����P�E��H�P��]� �����������������������U���D���3ŉE�VW�M̍E�P�M�"���M̃����P�Q�P�Q�@�A�M�Q�M�W���}̃��   ���_^�M�3��IC����]� ��������������������������������������U���D���3ŉE�VW�M̍E�P�M��!���M̃����P�Q�P�Q�@�A�M�Q�M�W���}̃��   ���_^�M�3��B����]� ��������������������������������������U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��j�h��d�    PQ��   ���3ŉE�SVWP�E�d�    �e��M��M��W���E��E�P�M��U���M��A    �U��B    �E��@    �E�    �M��t	�E��a�	�U��B�E��M�Q�M�U����p�����p���Rj �E�P�_/������x����M���x����Q�M�l���E��E�Pj �M�Q�!������|����U���|����B�M�(����t����M�Qj ��t���R�� �����E��E��M��H��M���B��j j ��T������E�������E������U��t0�E�Pj j.��<�����M�f�A�U�Rj j,��<�����M�f�A���,�   �u����U�Rj �M��vS���M�d�    Y_^[�M�3��5@����]� ������������������������������������������������������������������������������������������������������������������U��j�h��d�    PQ��   ���3ŉE�SVWP�E�d�    �e��M��M�U���E��E�P�M�S���M��A    �U��B    �E��@    �E�    �M��t	�E��a�	�U��B�E��M�Q�M�bS����p�����p���Rj �E�P�/-������x����M���x����Q�M��i���E��E�Pj �M�Q�$c������|����U���|����B�M�&����t����M�Qj ��t���R��b�����E��E��M��H��M��\��j j �R������E�������E������U��t0�E�Pj j.�n�����M�f�A�U�Rj j,��m�����M�f�A���,�   �u����U�Rj �M���!���M�d�    Y_^[�M�3��>����]� ������������������������������������������������������������������������������������������������������������������U��j�h �d�    PQ��SVW���3�P�E�d�    �e��M�E��@    �M��A    �U��B    �E�    �EPj �M��~I���M�h���E�M�U�Q��M���]��j j �;Q���x��E�������E������M�d�    Y_^[��]� ���������������������������������������������U��j�hP�d�    PQ��SVW���3�P�E�d�    �e��M�E��@    �M��A    �U��B    �E�    �EPj �M��=���M��g���E�M�U�Q��M��`,��j j �[P���X��E�������E������M�d�    Y_^[��]� ���������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M�E�P�M�D���E��M��M��E�    �U�R�M����(���E������M���c���M�d�    Y��]� �����������������������������U��j�h��d�    P�����3�P�E�d�    �M�E�P�M�
D���E��M��M��E�    �U�R�M���>(���E������M��]c���M�d�    Y��]� �����������������������������U��Q�M��} t#�M���.��9Er�M���.���M��Q�P;Ew2������]� ������������������U��Q�M��} t#�M��FK��9Er�M��9K���M��Q�P;Ew2������]� ������������������U��j�h �d�    P��   ���3ŉE�P�E�d�    h�  hx��EP�'�����}$ v�M ���+t�E ���-u	�E�   ��E�    �U��U��M��_��%   =   u@�E���;E$w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M��U�R�M��=����|�����|�����t����E�    ��t���Q��I�����E��E������M����j �U$R�M�����E�   j �M��-��P�E E$P�   k� U R�M��X���E�P�M�}=����x�����x����M��E��U�R�C�����E��E��M��0���E�P�M���9���E�j �M��"���E��M����tz�E����~p�M��4P��f�E��U����tY�M����~O�E���U$+U�;�s?�E���U$+щU$�E�Pj�M$Q�M��L���   �� �E����~	�U����U�뜍M���c���E$�M�\C���E��U��}� |%�}� v�M�@C��;E$v�M�3C��+E$�E���E�    �E��E��M��]��%�  �E��}�@ty�}�   tp�M�Q�UR�EP�MQ��T���R�EP��d������P�M�U�E�    �E�Pj �M���+��P�MQ�UR��l���P�MQ�WB������@�U�E�   �}�   um�M�Qj �M��+��P�UR�EP��D���Q�UR�B������P�M�U�E�P�MQ�UR�EP��\���Q�UR�d������P�M�U�E�    �5�E�Pj �M��6+��P�MQ�UR��L���P�MQ�A������@�U�E�M$+M�Q�U�R�M���*��P�EP�MQ��d���R�EP�mA������P�M�Uj j �M�'���E�P�MQ�UR�EP�MQ�UR�mc�����E��M��$%���E������M��-&���E�M�d�    Y�M�3���5����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h`�d�    P��   ���3ŉE�P�E�d�    h�  hx��EP�^�����}$ v�M ���+t�E ���-u	�E�   ��E�    �U��U��M�zZ��%   =   u@�E���;E$w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M��U�R�M�8����|�����|�����t����E�    ��t���Q�������E��E������M��E��j �U$R�M��V���E�   j �M��=��P�E E$P�   k� U R�M��(%���E�P�M�8����x�����x����M��E��U�R�i�����E��E��M������E�P�M��,���E�j �M��T���E��M����tz�E����~p�M�����f�E��U����tY�M����~O�E���U$+U�;�s?�E���U$+щU$�E�Pj�M$Q�M�����   �� �E����~	�U����U�뜍M��X���E$�M��=���E��U��}� |%�}� v�M��=��;E$v�M��=��+E$�E���E�    �E��E��M�xX��%�  �E��}�@ty�}�   tp�M�Q�UR�EP�MQ��T���R�EP��O������P�M�U�E�    �E�Pj �M���;��P�MQ�UR��l���P�MQ�;������@�U�E�   �}�   um�M�Qj �M��;��P�UR�EP��D���Q�UR��:������P�M�U�E�P�MQ�UR�EP��\���Q�UR�O������P�M�U�E�    �5�E�Pj �M��H;��P�MQ�UR��L���P�MQ�g:������@�U�E�M$+M�Q�U�R�M��;��P�EP�MQ��d���R�EP�-:������P�M�Uj j �M�+"���E�P�MQ�UR�EP�MQ�UR�cN�����E��M������E������M��==���E�M�d�    Y�M�3��d0����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P���   ���3�P�E�d�    j j �9!�����   ������#Uu�   �} um�pD���E�jUh��E�PjD�������E��E�    �}� tj �MQ�M���P���E���E�    �U�U��E���������\��P�E�P�M�Y'��� ����C��P�MQ�N?����P�M�7'��j j ��=�����   ������#Uu�   �} uy�C����P���jVh���P���Pj�9�����E��E�   �}� tj �MQ�M��%S���E���E�    �U���x����E�����������P��x���P�M�&��� ������P�MQ�U,����P�M�w&��j j �$�����   ������#Uu�   �} uy��B����8���jWh���8���Pj�y�����E��E�   �}� tj �MQ�M��
]���E���E�    �U؉�p����E������������P��p���P�M��%��� �������P�MQ�$����P�M�%��j j �Y%�����   ������#Uu�   �} u{�<B����H���jXh���H���Pj������E��E�   �}� tj j �MQ�M��$+���E���E�    �UЉ�h����E�����������P��h���P�M�%��� ������P�MQ�]7����P�M��$��j j �K/�����   ������#Uu�   �} uy�zA����(���jYh���(���Pj�������E��E�   �}� tj �MQ�M��D���E���E�    �Uȉ�`����E���������]��P��`���P�M�W$��� ����A��P�MQ��:����P�M�5$��j j �J�����   ������#Uu�   �} uy�@����@���jZh���@���Pj�7�����E��E�   �}� tj �MQ�M��X%���E���E�    �U���X����E�����������P��X���P�M�#��� ������P�MQ�DG����P�M�u#��j j �:�����   ������#Uu�   �} us��?����0���j[h���0���Pj�w�����E��E�   �}� tj �MQ�M���A���E���E�    �U�U��E������������P�E�P�M��"��� �������P�MQ�X����P�M�"��j j ��1�����   ������#Uu�   �} uy�@?����|���j\h���|���Pj������E��E�   �}� tj �MQ�M������E���E�    �U܉�t����E���������#��P��t���P�M�"��� ������P�MQ�5����P�M��!��j j �C�����   ������#Uu�   �} u{�>����l���j]h���l���PjX�������E��E�   �}� tj j �MQ�M��/V���E���E�    �Ủ�d����E���������a��P��d���P�M�[!��� ����E��P�MQ�-M����P�M�9!��j j �kY�����   ������#Uu�   �} u{�=����\���j^h���\���PjX�;�����E��E�	   �}� tj j �MQ�M��F���E���E�    �U���T����E�����������P��T���P�M� ��� ������P�MQ��'����P�M�w ��j j ������   ������#Uu�   �} uy��<����L���j_h���L���PjD�y�����E��E�
   �}� tj �MQ�M��-���E���E�    �U���D����E������������P��D���P�M����� �������P�MQ�����P�M���j j �������   ������#Uu�   �} uy�<<����<���j`h���<���Pj������E��E�   �}� tj �MQ�M��/?���E���E�    �U���4����E�����������P��4���P�M���� ������P�MQ�6A����P�M����j j �K&�����   ������#Uu�   �} uy�|;����,���jbh���,���Pj4�������E��E�   �}� tj �MQ�M��rJ���E���E�    �U���$����E���������_��P��$���P�M�Y��� ����C��P�MQ������P�M�7���M�d�    Y��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P���   ���3�P�E�d�    j j �������   ������#Uu�   �} um� 8���E�j-h��E�PjD������E��E�    �}� tj �MQ�M�����E���E�    �U�U��E������������P�E�P�M����� �������P�MQ�F����P�M����j j ��@�����   ������#Uu�   �} uy�L7����P���j.h���P���Pj�������E��E�   �}� tj �MQ�M������E���E�    �U���x����E���������/��P��x���P�M�)��� ������P�MQ�����P�M���j j �������   ������#Uu�   �} uy�6����8���j/h���8���Pj�	�����E��E�   �}� tj �MQ�M�������E���E�    �U؉�p����E���������o
��P��p���P�M�i��� ����S
��P�MQ�Z?����P�M�G��j j � �����   ������#Uu�   �} u{��5����H���j0h���H���Pj�I�����E��E�   �}� tj j �MQ�M������E���E�    �UЉ�h����E���������	��P��h���P�M���� ����	��P�MQ�������P�M���j j �.�����   ������#Uu�   �} uy�
5����(���j1h���(���Pj������E��E�   �}� tj �MQ�M��K���E���E�    �Uȉ�`����E������������P��`���P�M����� �������P�MQ�J����P�M����j j �5!�����   ������#Uu�   �} uy�J4����@���j2h���@���Pj�������E��E�   �}� tj �MQ�M�����E���E�    �U���X����E���������-��P��X���P�M�'��� ������P�MQ�� ����P�M���j j �2������   ������#Uu�   �} us�3����0���j3h���0���Pj������E��E�   �}� tj �MQ�M���/���E���E�    �U�U��E���������p��P�E�P�M�m��� ����W��P�MQ�a����P�M�K��j j �5������   ������#Uu�   �} uy��2����|���j4h���|���Pj�M�����E��E�   �}� tj �MQ�M��g���E���E�    �U܉�t����E�����������P��t���P�M���� ������P�MQ�������P�M���j j ������   ������#Uu�   �} u{�2����l���j5h���l���PjX������E��E�   �}� tj j �MQ�M��>>���E���E�    �Ủ�d����E������������P��d���P�M����� �������P�MQ�����P�M����j j �`�����   ������#Uu�   �} u{�N1����\���j6h���\���PjX�������E��E�	   �}� tj j �MQ�M���>���E���E�    �U���T����E���������/��P��T���P�M�)��� ������P�MQ��>����P�M���j j � �����   ������#Uu�   �} uy�0����L���j7h���L���PjD�	�����E��E�
   �}� tj �MQ�M��'���E���E�    �U���D����E���������o��P��D���P�M�i��� ����S��P�MQ��J����P�M�G��j j �S5�����   ������#Uu�   �} uy��/����<���j8h���<���Pj�I�����E��E�   �}� tj �MQ�M��s����E���E�    �U���4����E�����������P��4���P�M���� ������P�MQ�&����P�M���j j �������   ������#Uu�   �} uy�/����,���j:h���,���Pj4�
�����E��E�   �}� tj �MQ�M���D���E���E�    �U���$����E������������P��$���P�M����� �������P�MQ�
����P�M�����M�d�    Y��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EP�?!�������E�jAh`���+��P3ɋE��   �������Q�n������E�E�E��M�Q�UR�E�P� 5�����E���]����������������������������U����M��E��H(��u,�}w&�}w �}wkU�E��kU(��x��E���E�Ȧ�M��M�j�U�Rj�EP��������]� �������������������������U����M��E��H(��u,�}w&�}w �}wkU�E��kU(��x��E���E�Ȧ�M��M�j�U�Rj�EP�J������]� �������������������������U����M��E��xr�M��QR�!�����E��	�E����E��E���]���������������������������U����M��E��xr�M��QR�������E��	�E����E��E���]���������������������������U����M��E��xr�M��QR������E��	�E����E��E���]���������������������������U����M��E��xr�M��QR�Y�����E��	�E����E��E���]���������������������������U��j�hp�d�    P�����3�P�E�d�    �E�   �} u	�E�    ��EP�M�}8���E��M��M��E� �M�����E������M�����E�M�d�    Y��]������������������������������������U��j�h��d�    P�����3�P�E�d�    �E�   �} u	�E�    ��EP�M�[2���E��M��M��E� �M�l����E������M�]����E�M�d�    Y��]������������������������������������U����M�E�8 t.�M�	�	��f�E���%��f�E��U�R�E�P�������ȅ�t�U��    ��E�P�O-�����M�f�A�U��B�E�f�@��]����������������������������������U����M�E�8 t.�M�	����f�E��&;��f�E��U�R�E�P��5�����ȅ�t�U��    ��E�P������M�f�A�U��B�E�f�@��]����������������������������������U����M��E��H �9 t�U��B0��M���E�    �E����]�����������������U����M��E��H �9 t�U��B0��M���E�    �E����]�����������������U����M��E��H0����E��H0��U��B ��M��U��B ����U��B ��E���]��������������������������������U����M��E��H0����E��H0��U��B ��M��U��B ����U��B ��E���]��������������������������������U��j�h��d�    P���3�P�E�d�    �E�    ��E ���E �M�08���M� '���}  v �M����f���R�M������ �����E�M��U�P�E������M������E�M�d�    Y��]����������������������������������������U��j�h�d�    P���3�P�E�d�    �E�    ��E ���E �M�����M�-���}  v �M�-��f���R�M������������E�M��U�P�E������M�����E�M�d�    Y��]����������������������������������������U����E���E�M��6���M���M�} v�U�P�M�7��������ȋM�U��E�A�E]���������������������������������U����E���E�M�����M���M�} v�U�P�M����������ȋM�U��E�A�E]���������������������������������U��j�h��d�    P��  ���3ŉE�P�E�d�    ��X����E�    h  h��EP�������M��tK������R�M����������������������E�������Q�]������8����E� �����������I��t���R�M������������������|����E���|���Q�1������8����E� ��t����h����U�R��8���� ���E���8���������������� }������؉����������������������@����M$�S8��;�@���w(�E@P�M$�>8����@���+ȃ�Qj �M$�6 ����   �M��T��������   �M��@���� ����   ��8����7��f������M�������0����M$��7��+�@�����(�����0������tx��0������~k��0����;�(���sZ��0������(���+�(��������Qj��(���R�M$�z���   �� ��0������~��0�������0����z����M��2:���E��M ��tH��`���R��8����d���� �� ����M�Q��8���������x�����x���R�M������M��L����L��H���P��8���������� �����H���R��8�������������������P�M��4�����H���������M��9���E��M��0����t2��d���Q��8����&��������������R�M��������d�������ƅ?��� ǅD���    ǅ4���    ���4�������4�����4����  ��4����� �����,�����,����� ��,�����,���X��   ��,������B�$��B�M���5���D�����D����   �M��5���D�����D����   ��@��� vǅ���   �
ǅ���    �M$�y5��;�@���w�M$�i5����@���+ȃ�������
ǅ���    �M$�D5�����������D�����D������D�������D�����4���tƅ?���������M��������������������� |1	������ v&�M�o��;�D���v�M�_��+�D���������
ǅ���    �������D����M��.��%�  ����������@tO�����   u��?�����u8��D���R�EP�MQ�UR������P��������P�M�UǅD���    ǅ4���    ���4�������4�����4����  ��4����� �����$�����$����� ��$�����$���X��  ��$�����4C�$�C�M���3��P�����P�M�������������������������E����̉�@���������R�5����8����EP�MQ������R�7������������������P�M�U�E�������W����5  �M��63������   j��$���P�M��4����������������������E����̉�0���������R�5����L����EP�MQ������R��6������������������P�M�U�E���$���������  ��@��� ��   �M$�2��P�����P�M$�����������������������E����̉�P���������R�r4����p����EP�MQ������R�e6������������������P�M�U�E�������'����  �M$�2��;�@����	  �E@Pj �M�J������������X����8����7����Qj �M�#�����������1���M$�1����@���+�R�E@P�MQ�UR��|���P���������P�M�U�M$�v1��P������P�M$�}����������������������E�	���̉�d���������R�U3����<����EP�MQ��l���R�H5������������������P�M�U�E��������
����y  �M$��0��+�@���P������P�M$������������������������E�
���̉�\���������R��2����D����EP�MQ��t���R�4������������������P�M�U�E��������w�����8����5����Pj �M�������4���������@���Q��@���R������P������Q�M$�����������������������E��������/���������������������E����̉�T���������R��1����4����EP�MQ������R��3������������������P�M�U�E������������E������������mj�EP�MQ�UR������P��������P�M�U�����   u8��D���P�MQ�UR�EP������Q�u�������@�U�EǅD���    ������M���.������   �M���.����Pj�� ���Q������R�M�������������������� ����E��� ���������������������������E����̉�l���������R�0����h����EP�MQ������R�2������������������P�M�U�E��� ����R����E��������C���j j �M������D���P�MQ�UR�EP�MQ�Z������E��M��[����E��M��O����E� �M��+����E������M$�4����E�M�d�    Y�M�3�������]�< 0;�:�:�:?;O; �I �@�<=�=AQA ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��  ���3ŉE�P�E�d�    ��X����E�    h  h��EP�'�����M��tK������R�M����������������������E�������Q�� ������8����E� �����������I��t���R�M������������������|����E���|���Q���������8����E� ��t����h����U�R��8���������E���8�����-������������ }������؉����������������������@����M$�"��;�@���w(�E@P�M$�"����@���+ȃ�Qj �M$�D�����   �M��T��������   �M��@���� ����   ��8����!��f������M�������0����M$�"��+�@�����(�����0������tx��0������~k��0����;�(���sZ��0������(���+�(��������Qj��(���R�M$�����   �� ��0������~��0�������0����z����M��W
���E��M ��tH��`���R��8������� �� ����M�Q��8���������x�����x���R�M������M�����L��H���P��8���������� �����H���R��8������������������P�M�������H����n���M��	���E��M�� ����t2��d���Q��8����|���������������R�M��n�����d����#��ƅ?��� ǅD���    ǅ4���    ���4�������4�����4����  ��4����� �����,�����,����� ��,�����,���X��   ��,������R�$��R�M�� ���D�����D����   �M������D�����D����   ��@��� vǅ���   �
ǅ���    �M$����;�@���w�M$�����@���+ȃ�������
ǅ���    �M$������������D�����D������D�������D�����4���tƅ?���������M��������������������� |1	������ v&�M�o��;�D���v�M�_��+�D���������
ǅ���    �������D����M����%�  ����������@tO�����   u��?�����u8��D���R�EP�MQ�UR������P��������P�M�UǅD���    ǅ4���    ���4�������4�����4����  ��4����� �����$�����$����� ��$�����$���X��  ��$�����4S�$�S�M��
��P�����P�M��T���������������������E����̉�@���������R������8����EP�MQ������R�������������������P�M�U�E������������5  �M��}������   j��$���P�M�����������������������E����̉�0���������R������L����EP�MQ������R�"������������������P�M�U�E���$����,����  ��@��� ��   �M$����P�����P�M$�$���������������������E����̉�P���������R������p����EP�MQ������R�������������������P�M�U�E�����������  �M$�M��;�@����	  �E@Pj �M�R�����������������8����������Qj �M�+����������������M$������@���+�R�E@P�MQ�UR��|���P�B�������P�M�U�M$���P������P�M$����������������������E�	���̉�d���������R�e�����<����EP�MQ��l���R�k������������������P�M�U�E��������u����y  �M$�0��+�@���P������P�M$�t���������������������E�
���̉�\���������R�������D����EP�MQ��t���R��������������������P�M�U�E��������������8����k�����Pj �M�������{������> ����@���Q��@���R������P������Q�M$�����������������������E��������o����������������������E����̉�T���������R�������4����EP�MQ������R��������������������P�M�U�E������������E�������������mj�EP�MQ�UR������P��������P�M�U�����   u8��D���P�MQ�UR�EP������Q���������@�U�EǅD���    ������M��C������   �M��2����Pj�� ���Q������R�M��p���������������� ����E��� ����c���������������������E����̉�l���������R������h����EP�MQ������R�������������������P�M�U�E��� ��������E�����������j j �M������D���P�MQ�UR�EP�MQ�������E��M�������E��M������E� �M��+����E������M$�����E�M�d�    Y�M�3��������]�< 0K�J�J�J?KOK �I �P�LM�MQQQ ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E���E�M�����} v�MQ�M�b�����������ӋU�E��M�J�E]����������������������������U����E���E�M�����} v�MQ�M�I����������ӋU�E��M�J�E]����������������������������U����E���E�M�6���} v�MQ�M�������%����ӋU�E��M�J�E]����������������������������U����E���E�M������} v�MQ�M�������L����ӋU�E��M�J�E]����������������������������U��Q�M��E��HQ��������U��BP��������M��QR��������E��HQ���������]��������������������������U��Q�M��E��HQ�������U��BP�������M��QR�r������E��HQ�c�������]��������������������������U����M��E��u�s�M��yrj�U��B�E�M���Q�U�R�M��������F���} v �EP�M�Q�m�����P�U���R�������E��H��Q�U�R�E�P�M��l����������M��A   �UR�M��������]� ����������������������������������������������U����M��E��u�s�M��yrj�U��B�E�M���Q�U�R�M����������	���} v �EP�M�Q�������P�U���R�������E��H��Q�U�R�E�P�M������������M��A   �UR�M��������]� ����������������������������������������������U��Q�M��E��HQ�������U��BP�������M��QR�r�������]�������������������������U��Q�M��E��HQ�@������U��BP�1������M��QR�"�������]�������������������������U��Q�M��E��HQ��������U��BP��������M��QR���������]�������������������������U��Q�M��E��HQ�������U��BP�������M��QR��������]�������������������������U����M��1	���E��}� t�E�P�M����"����M�Q�������M�������Ѕ�u�M��������E���E�x��E��]�������������������������������U����M������E��}� t�E�P�M��������M�Q�I�����M����)���Ѕ�u�M����4����E���E�H��E��]�������������������������������U����M��E�    ����P�M�����E����E��E��]� ����������������U��Q�M�hm�[����]������������U��Q�M�hm�;����]������������U��Q�M�h m�������]������������U��Q�M�h m������]������������U��Q�M��EP�M�������]� �������U��Q�M��EP�M��������]� �������U��Q�M�j �EP�	������]� ���������������������U��Q�M�j �EP���������]� ���������������������U��Q�M��P�Pj �MQ�M������]� ���������������U����M��M����;Es�M��;����M����+E�E��E�;Es�M��M�U��P�+B;Ew�M������} vZ�M��QU�U�j �E�P�M������ȅ�t9�UR�M�����M�HR�M������M��Q�PP��������M�Q�M��a����E���]� �����������������������������������������������������U����M��E��P�+H;Mw�M�����} vE�U��BE�E�j �M�Q�M��
���Ѕ�t$�EP�MQ�U��BP�M��P����M�Q�M������E���]� ������������������������������������������U��Q�M����Pj �MQ�M�������]� ���������������U����M��M�`
��;Es�M������M�K
��+E�E��E�;Es�M��M�U����+B;Ew�M��q���} vZ�M��QU�U�j �E�P�M������ȅ�t9�UR�M�R����M�HR�M������M��Q�PP� ������M�Q�M��p����E���]� �����������������������������������������������������U����M��E����+H;Mw�M�����} vE�U��BE�E�j �M�Q�M�������Ѕ�t$�EP�MQ�U��BP�M��p����M�Q�M�������E���]� ������������������������������������������U����M��E�;Eu�a�M�Q�M�g���P�U�R�M��Z���P�����������t�M�yr�UR�M������!j j�M������EP������P�M������E���]� �����������������������������������U��Q�M��P�Pj �MQ�M������]� ���������������U����M��M���;Es�M������M���+E�E��E;E�s�M�M��U�;Uu�EE�P�M��-����MQj �M��v����Ej �U�R�M��������t0�M�Q�M�v����U�PP�M�����P��������M�Q�M��M����E���]� �������������������������������������������������U��Q�M��E;P�u�M�����j �MQ�M�����Ѕ�t�EP�MQj �M��_����UR�M�������E���]� �������������������������U��Q�M�h�  h ��EP�u������MQ������P�UR�M��	�����]� ��������������������U��Q�M��} th  h ��EP�������MQ�M��d���Ѕ�t"�EP�M��M����M+���Q�U�R�M�� ���=j �EP�M��
���ȅ�t%�UR�EP�M�����P�:������MQ�M�������E���]� �����������������������������������������������������U����M��E�;Eu�a�M�Q�M����P�U�R�M�����P�� ��������t�M�yr�UR�M�������!j j�M�������EP蓿����P�M��S����E���]� �����������������������������������U��Q�M����Pj �MQ�M��\�����]� ���������������U����M��M����;Es�M��l����M���+E�E��E;E�s�M�M��U�;Uu�EE�P�M������MQj �M�菿���Ej �U�R�M��!�������t0�M�Q�M�����U�PP�M��
���P�l������M�Q�M�������E���]� �������������������������������������������������U��Q�M��E;��u�M��)��j �MQ�M������Ѕ�t�EP�MQj �M�������UR�M��T����E���]� �������������������������U��Q�M�h�  h ��EP�������MQ�:�����P�UR�M�������]� ��������������������U��Q�M��} th  h ��EP�7������MQ�M������Ѕ�t"�EP�M������M+���Q�U�R�M��Q����=j �EP�M������ȅ�t%�UR�EP�M��~���P��������MQ�M��P����E���]� �����������������������������������������������������U��EP�MQ�UR�������]�������U��E�Mf�f�]����������������U��EP�MQ�UR������]�������U��E�Mf�f�]����������������U��Q�M��E�P�M������P�M�/���E��]� �����������U��Q�M��E�P�M��h���P�M������E��]� �����������U��Q�M��M��Y�����]��������������U��Q�M��M�������]��������������U��Q�} u�E�E���MQ�UR�EP��������E��E���]�����������������U��Q�} u�E�E���MQ�UR�EP�������E��E���]�����������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M��EP�MQ�M���	����]� �������������������U��Q�M��EP�MQ�M�������]� �������������������U��Q�M��EP� 	������]� �������U��Q�M��EP��������]� �������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M�2���]����U��Q�M�2���]����U��Q�M���]� ���U��Q�M���]� ���U����M�j_hP��EP�MQ������j`hP��UR�EP�������M���Q�UR�EP�MQ�UR��������E��}� }	�E�������}� u	�E�    ��E�   �E��E�E��]� �����������������������������������U����M�j_hP��EP�MQ�������j`hP��UR�EP�������M���Q�UR�EP�MQ�UR�t�����E��}� }	�E�������}� u	�E�    ��E�   �E��E�E��]� �����������������������������������U����M��E�    �E��HQ�M�
����U����U��E��]� ���������������U����M��E�    �E��HQ�M�����U����U��E��]� ���������������U��Q�M��E��@��]����������������U��Q�M��E��@��]����������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M�3���]����U��Q�M�3���]����U����M��E�    �E��HQ�M誾���U����U��E��]� ���������������U����M��E�    �E��HQ�M�6����U����U��E��]� ���������������U��Q�M��E��@��]����������������U��Q�M��E��@��]����������������U����M��E�    �EP�M�y����M����M��E��]� ������������������U����M��E�    �EP�M�n����M����M��E��]� ������������������U��j�hH�d�    P��P���3ŉE�P�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M�������E�    �EP�MQ�v������Ѕ�t�E$����U$�
�M��
�����u�E$����U$�
�P�M�������E��E�    �E�Pj �M�Q�U�R��������]��E�;E�t�}� t�M$����E$���M(�E���U�E��M�J�E������M������E�M�d�    Y�M�3��V�����]�$ �����������������������������������������������������������������������������������U��j�h��d�    P��H���3ŉE�VP�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M������E�    �M������E��EP�MQ��������Ѕ�t�E$����U$�
�}� u�E$����U$�
�   �E�    �E�P�M(�����j �M��%������-u+�U��U��E�P�M(������   k�
f�L�f��U����U��	�E����E��M�;M�s(�U�R�M��Ӻ���0�E�P�M(����f��ux���f��ǋU�E��M�J�E������M�������E�M�d�    Y^�M�3�������]�$ ����������������������������������������������������������������������������������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M�������E�    �EP�MQ�^������Ѕ�t�E$����U$�
�M��������u�E$����U$�
�P�M��ɹ���E��E�    �E�Pj �M�Q�U�R��������]��E�;E�t�}� t�M$����E$���M(�E���U�E��M�J�E������M��w����E�M�d�    Y�M�3��&�����]�$ �����������������������������������������������������������������������������������U��j�h�d�    P��H���3ŉE�VP�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M��c����E�    �M������E��EP�MQ�������Ѕ�t�E$����U$�
�}� u�E$����U$�
�   �E�    �E�P�M(�4���j �M���������-u+�U��U��E�P�M(�����   k�
f�L�f��U����U��	�E����E��M�;M�s(�U�R�M�裷���0�E�P�M(�����f��ux���f��ǋU�E��M�J�E������M��ý���E�M�d�    Y^�M�3��q�����]�$ ����������������������������������������������������������������������������������������������U��j�hH�d�    P��P���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP��������E�    �M�Q�M�q����E��U��U��E�    �E�P�M�����P�MQ�UR�E�P�M�Q�X������E��E������M������   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R�������E̍EP�MQ�������Ѕ�t�E ����U �
�E�;E�t�}� u	�}���  v�M ����E ��,�   k� �DЃ�-u
3�+M̉M���ỦUċE$f�M�f��U�E��M�J�E�M�d�    Y�M�3�������]�  ������������������������������������������������������������������������������������������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP��������E�    �M�Q�M�����E��U��U��E�    �E�P�M�����P�MQ�UR�E�P�M�Q�h������E��E������M������   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R�������E̍EP�MQ�������Ѕ�t�E ����U �
�E�;E�t�}� u�}��v�M ����E ��*�   k� �DЃ�-u
3�+M̉M���ỦUċE$�Mĉ�U�E��M�J�E�M�d�    Y�M�3�������]�  �����������������������������������������������������������������������������������������������������������U��j�h��d�    P��@���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP��������E�    �M�Q�U�R�M�����E��E��E��E�    �M�Q�M�����P�UR�EP�M�Q�U�R�t�����P�E�P�M�Q�-������E��E������M������UR�EP��������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3�������]�  �������������������������������������������������������������������������������U��j�h�d�    P��@���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP�f������E�    �M�Q�U�R�M�����E��E��E��E�    �M�Q�M�u���P�UR�EP�M�Q�U�R�������P�E�P�M�Q�a������E��E������M�薥���UR�EP�M������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3�������]�  �������������������������������������������������������������������������������U���T���3ŉE��M�h)  hx��EP�MQ�UR�EP��������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q�	�����P�U�R�E�P��������]��}� t�M���QQ�E��$�������]��UR�EP��������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��/�����]�  ����������������������������������������������������������������������������U���X���3ŉE��M�hA  hx��EP�MQ�UR�EP�������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q������P�U�R�E�P�`������]��}� t�M���Q���E��$趡�����]��UR�EP�������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��������]�  ��������������������������������������������������������������������������U���X���3ŉE��M�hY  hx��EP�MQ�UR�EP�^������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q�i�����P�U�R�E�P�[������]��}� t�M���Q���E��$�U������]��UR�EP�M������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3�������]�  ��������������������������������������������������������������������������U��j�hH�d�    P��P���3ŉE�P�E�d�    �M�hq  hx��EP�MQ�UR�EP��������E�    �M�Q�M�����E��U��U��E�    �E�Ph   �MQ�UR�E�P�M�Q茽�����E��E������M��?����   ��t"�E�P�M�Q�U�R�E�P�������3ɉE��M���U�R�E�P�M�Q�U�R�������E��U��E��E��M��M��UR�EP�������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E��M$��U�E��M�J�E�M�d�    Y�M�3��������]�  ���������������������������������������������������������������������������������������������������U��j�h��d�    P��D���3ŉE�P�E�d�    �M�h   hx��EP�MQ�UR�EP�&������E�    �M�Q�U�R�M������E��E��E��E�    �M�Q�M�5���P�UR�EP�M�Q�U�R贻����P�E�P�M�Q�+������E��U��E������M��S����UR�EP�
������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3��9�����]�  ��������������������������������������������������������������������������������������U��j�h��d�    P��D���3ŉE�P�E�d�    �M�h  hx��EP�MQ�UR�EP�������E�    �M�Q�U�R�M�=����E��E��E��E�    �M�Q�M����P�UR�EP�M�Q�U�R�$�����P�E�P�M�Q�t������E��U��E������M��Ü���UR�EP�z������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3�詾����]�  ��������������������������������������������������������������������������������������U��j�h1�d�    P��   ���3ŉE�P�E�d�    ��L���h�  hx��EP�MQ�UR�EP� �����ǅx��������M�0���% @  �'  ��H���Q�M������\�����\�����P����E�    ��P���P���������p����E�������H����3���j j�M��,����E�   ��|���Q��p����յ����@�����@�����8����E���8���P�M��<����E���|���膭��j �M������M�Q��p���蛢����d�����d�����<����E���<���P�M�������E��M��<����M������Pj�MQ�UR虿������x����E������M������   ǅh���    ��h���P��`���Q�M�Z�����T�����T�����D����E�   ��D���P�M����P�MQ�UR�E�P��L���Q�2�����P��X���R�E�P��������l����E�������`����˙���M�9�X���t��h��� u��l���w��l�����x����EP�MQ�Y������Ѕ�t�E ����U �
��x��� }�E ����U �
�*��x��� tǅt���   �
ǅt���    �E$��t�����U�E��M�J�E�M�d�    Y�M�3��q�����]�  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hx�d�    P��P���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP��������E�    �M�Q�M�����E��U��U��E�    �E�P�M�y���P�MQ�UR�E�P�M�Q�r������E��E������M�諗���   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R�&������E̍EP�MQ�9������Ѕ�t�E ����U �
�E�;E�t�}� u	�}���  v�M ����E ��,�   k� �DЃ�-u
3�+M̉M���ỦUċE$f�M�f��U�E��M�J�E�M�d�    Y�M�3��)�����]�  ������������������������������������������������������������������������������������������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP��������E�    �M�Q�M�!����E��U��U��E�    �E�P�M����P�MQ�UR�E�P�M�Q肻�����E��E������M�軕���   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R�6������E̍EP�MQ�I������Ѕ�t�E ����U �
�E�;E�t�}� u�}��v�M ����E ��*�   k� �DЃ�-u
3�+M̉M���ỦUċE$�Mĉ�U�E��M�J�E�M�d�    Y�M�3��>�����]�  �����������������������������������������������������������������������������������������������������������U��j�h��d�    P��@���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP�������E�    �M�Q�U�R�M�-����E��E��E��E�    �M�Q�M����P�UR�EP�M�Q�U�R莹����P�E�P�M�Q�͹�����E��E������M�趓���UR�EP腞�����ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3�袵����]�  �������������������������������������������������������������������������������U��j�h8�d�    P��@���3ŉE�P�E�d�    �M�h�  hx��EP�MQ�UR�EP�������E�    �M�Q�U�R�M譹���E��E��E��E�    �M�Q�M����P�UR�EP�M�Q�U�R������P�E�P�M�Q�������E��E������M��6����UR�EP�������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3��"�����]�  �������������������������������������������������������������������������������U���T���3ŉE��M�h)  hx��EP�MQ�UR�EP�%������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q�%�����P�U�R�E�P�i������]��}� t�M���QQ�E��$�[������]��UR�EP觛�����ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��ϲ����]�  ����������������������������������������������������������������������������U���X���3ŉE��M�hA  hx��EP�MQ�UR�EP��������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q�չ����P�U�R�E�P� ������]��}� t�M���Q���E��$�V������]��UR�EP�U������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��}�����]�  ��������������������������������������������������������������������������U���X���3ŉE��M�hY  hx��EP�MQ�UR�EP�������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q腸����P�U�R�E�P��������]��}� t�M���Q���E��$��������]��UR�EP�������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��-�����]�  ��������������������������������������������������������������������������U��j�hx�d�    P��P���3ŉE�P�E�d�    �M�hq  hx��EP�MQ�UR�EP�������E�    �M�Q�M�A����E��U��U��E�    �E�Ph   �MQ�UR�E�P�M�Q覲�����E��E������M��ߌ���   ��t"�E�P�M�Q�U�R�E�P�w�����3ɉE��M���U�R�E�P�M�Q�U�R�8������E��U��E��E��M��M��UR�EP�Y������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E��M$��U�E��M�J�E�M�d�    Y�M�3��v�����]�  ���������������������������������������������������������������������������������������������������U��j�h��d�    P��D���3ŉE�P�E�d�    �M�h   hx��EP�MQ�UR�EP�M������E�    �M�Q�U�R�M�m����E��E��E��E�    �M�Q�M�����P�UR�EP�M�Q�U�R�ΰ����P�E�P�M�Q�˻�����E��U��E������M������UR�EP������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3��٬����]�  ��������������������������������������������������������������������������������������U��j�h��d�    P��D���3ŉE�P�E�d�    �M�h  hx��EP�MQ�UR�EP�������E�    �M�Q�U�R�M�ݰ���E��E��E��E�    �M�Q�M�E���P�UR�EP�M�Q�U�R�>�����P�E�P�M�Q�������E��U��E������M��c����UR�EP�2������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3��I�����]�  ��������������������������������������������������������������������������������������U��j�ha d�    P��   ���3ŉE�P�E�d�    ��L���h�  hx��EP�MQ�UR�EP�'�����ǅx��������M�����% @  �'  ��H���Q�M�2�����\�����\�����P����E�    ��P���P�u�������p����E�������H����Ӈ��j j�M������E�   ��|���Q��p����=�����@�����@�����8����E���8���P�M��I����E���|���薶��j �M��@����M�Q��p����n�����d�����d�����<����E���<���P�M�������E��M��L����M��Ҿ��Pj�MQ�UR�;�������x����E������M������   ǅh���    ��h���P��`���Q�M�������T�����T�����D����E�   ��D���P�M�V���P�MQ�UR�E�P��L���Q�L�����P��X���R�E�P�<�������l����E�������`����k����M�9�X���t��h��� u��l���w��l�����x����EP�MQ�������Ѕ�t�E ����U �
��x��� }�E ����U �
�*��x��� tǅt���   �
ǅt���    �E$��t�����U�E��M�J�E�M�d�    Y�M�3�������]�  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h� d�    P��p���3�P�E�d�    �M��E�P�M�ݫ���E܋M܉M��E�    �U�R�ѷ�����E��E������M�萄���E�    �E(�E�M��A�M�}�8�K  �U������$�D��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��Y�����P�M�U�  �E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�蹖����@�U�E��  h(��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��i�����P�M�U�  �E�P�M�Qjcj �UR�EP�M�Q�Ѝ�����U �M ��U ���ukM�d��l  �U$�J�Q  �E�P�M$��Qjj�UR�EP�M�Q脍�����U �M ��  hD��U$R�E P�MQ�UR�EP�MQ�UR�E�P�M�������P�M�U��  �E�P�M$��Qjj �UR�EP�M�Q�������U �M ��  �U�R�E$��Pjj �MQ�UR�E�P�������M �U ��~  �E�P�M$��Qhn  j�UR�EP�M�Q讌�����U �M ��I  �U�R�E�Pjj�MQ�UR�E�P�������M �U ��E ���u�U���E$�P�  �M�Q�U$��Rj;j �EP�MQ�U�R�7������M �U ���  hT��E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��d�����@�U�E�  hX�j �MQ�UR�ސ�����E�}� }�E ����U �
�kE��M$A�U$�B�Q  hh��E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��������@�U�E�  h|��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�������P�M�U��  �E�P�M$Qj;j �UR�EP�M�Q�������U �M ��  h���U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��:�����P�M�U�k  �E�P�M$��Qj5j �UR�EP�M�Q螊�����U �M ��9  �U�R�E$��Pjj �MQ�UR�E�P�l������M �U ��  �E�P�M$��Qj5j �UR�EP�M�Q�:������U �M ���   h���U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��g�����P�M�U�   �E�P�M�Qjcj �UR�EP�M�Q�Ή�����U �M ��U ���u �}�E}�M��d�M���U�U��E$�M��H�B�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��n�����P�M�U��E ����U �
�EP�MQ�Φ�����Ѕ�t�E ����U �
�E�M��U�P�E�M�d�    Y��]�( �I ���a�ܞ�K����$�S�������$���}���)�f���¡&�c�� 	
	 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h� d�    P��p���3�P�E�d�    �M��E�P�M�m����E܋M܉M��E�    �U�R��~�����E��E������M�� |���E�    �E(�E�M��A�M�}�8�K  �U�����$����M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��2~����P�M�U�  �E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�谟����@�U�E��  h(��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�������P�M�U�  �E�P�M�Qjcj �UR�EP�M�Q蓬�����U �M ��U ���ukM�d��l  �U$�J�Q  �E�P�M$��Qjj�UR�EP�M�Q�G������U �M ��  hD��U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��������P�M�U��  �E�P�M$��Qjj �UR�EP�M�Q�ث�����U �M ��  �U�R�E$��Pjj �MQ�UR�E�P覫�����M �U ��~  �E�P�M$��Qhn  j�UR�EP�M�Q�q������U �M ��I  �U�R�E�Pjj�MQ�UR�E�P�B������M �U ��E ���u�U���E$�P�  �M�Q�U$��Rj;j �EP�MQ�U�R��������M �U ���  hT��E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�胿����@�U�E�  hX�j �MQ�UR跼�����E�}� }�E ����U �
�kE��M$A�U$�B�Q  hh��E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�������@�U�E�  h|��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��ž����P�M�U��  �E�P�M$Qj;j �UR�EP�M�Q�Щ�����U �M ��  h���U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��Y�����P�M�U�k  �E�P�M$��Qj5j �UR�EP�M�Q�a������U �M ��9  �U�R�E$��Pjj �MQ�UR�E�P�/������M �U ��  �E�P�M$��Qj5j �UR�EP�M�Q��������U �M ���   h���U$R�E P�MQ�UR�EP�MQ�UR�E�P�M�膽����P�M�U�   �E�P�M�Qjcj �UR�EP�M�Q葨�����U �M ��U ���u �}�E}�M��d�M���U�U��E$�M��H�B�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M�蔙����P�M�U��E ����U �
�EP�MQ�v������Ѕ�t�E ����U �
�E�M��U�P�E�M�d�    Y��]�( �I $�\�ѦL�����g�W���é �d�)�����"���֨�2���Ӫ^� 	
	 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hd�    P��D���3�P�E�d�    �M�h  h���EP�MQ�UR�EP�)�����h  h���M$Q�M������U�R�M�Ś���E��E��E��E�    �M�Q蹦�����E��E������M��xs���M�蜫���E�}� u�E�   �UR�EP�������ȅ�t�  �M趏����Rj�M��+�������u?�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�躅����P�M�U�E�   �   �}�u>�E�P�M$��Qjj�UR�EP�M�Q��|�����U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P�|�����M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��{����@�U�E�MQ�UR�ؾ��������t'�M藎����QjH�M������Ѕ�t
�M������EP�MQ蚾�����Ѕ�t<j �M�W�����P�M������E��M��:t�U��,t	�E��/u�M詠���MQ�UR�G���������t'�M������QjH�M��{����Ѕ�t
�M�m����EP�MQ�$������Ѕ�t��   �M�Í����Pj�M��8����ȅ�uW�}�u�U ����M ��@�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M�貃����P�M�U�}�u�E�   �w�}�t�}�u>�E�P�M$��Qjj�UR�EP�M�Q��z�����U �M ��U$�B���M$�A�-�U�R�E$��Pjj�MQ�UR�E�P�z�����M �U ��EP�MQ�������Ѕ�t'�M�������PjH�M��6����ȅ�t
�M�(����UR�EP�ļ�����ȅ�t<j �M职����R�M������E��E��:t�M��,t	�U��/u�M�Ӟ���EP�MQ�q������Ѕ�t'�M�0�����PjH�M�襸���ȅ�t
�M藞���UR�EP�N������ȅ�t�U ����M ��  �M�������Rj�M��U�������uM�}�t�M ����E ��3�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��ρ����P�M�U�   �}�u>�E�P�M$��Qjj�UR�EP�M�Q�y�����U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P��x�����M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��w����@�U�E�MQ�UR����������t�M ����E ��M�U��E�A�E�M�d�    Y��]�  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h8d�    P��D���3�P�E�d�    �M�h  h���EP�MQ�UR�EP�0�����h  h���M$Q�ͺ�����U�R�M�E����E��E��E��E�    �M�Q�n�����E��E������M���k���M��m���E�}� u�E�   �UR�EP�v�����ȅ�t�  �M�1�����Rj�M��^�������u?�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�衏����P�M�U�E�   �   �}�u>�E�P�M$��Qjj�UR�EP�M�Q豜�����U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P�m������M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�蚍����@�U�E�MQ�UR����������t'�M������QjH�M��?����Ѕ�t
�M�����EP�MQ�ۇ�����Ѕ�t<j �M�Қ����P�M���o���E��M��:t�U��,t	�E��/u�M苯���MQ�UR與��������t'�M聚����QjH�M�讇���Ѕ�t
�M�O����EP�MQ�t�����Ѕ�t��   �M�>�����Pj�M��k����ȅ�uW�}�u�U ����M ��@�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M�虍����P�M�U�}�u�E�   �w�}�t�}�u>�E�P�M$��Qjj�UR�EP�M�Q蠚�����U �M ��U$�B���M$�A�-�U�R�E$��Pjj�MQ�UR�E�P�b������M �U ��EP�MQ�C������Ѕ�t'�M�<�����PjH�M��i����ȅ�t
�M�
����UR�EP�������ȅ�t<j �M�������R�M���m���E��E��:t�M��,t	�U��/u�M赭���EP�MQ貅�����Ѕ�t'�M諘����PjH�M��؅���ȅ�t
�M�y����UR�EP��r�����ȅ�t�U ����M ��  �M�[�����Rj�M�舅������uM�}�t�M ����E ��3�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�趋����P�M�U�   �}�u>�E�P�M$��Qjj�UR�EP�M�Q�͘�����U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P艘�����M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�趉����@�U�E�MQ�UR�q��������t�M ����E ��M�U��E�A�E�M�d�    Y��]�  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M�h}  h���EP�MQ�UR�EP�H�����h~  h���M$Q�l������U��BPj �MQ�UR�܉�����E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U����M�h}  h���EP�MQ�UR�EP������h~  h���M$Q謲�����U��BPj �MQ�UR�������E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U��j�hhd�    P�����3�P�E�d�    �M�h�   h���EP�MQ�UR�EP詯����h�   h���M$Q�ͱ�����U�R�M�E����E�E�E��E�    �M�Q�9������E��E������M���b���U�R�E$��Pjj �MQ�UR�E�P�m�����M �U ��E �8 uj �M�3����Q�M��ʁ���Ѓ�:t�E ����U �
�2�E�P�M$��Qj;j �UR�M�y���P�E�P�l�����M �U ��E �8 uj �M��~����Q�M��c����Ѓ�:t�E ����U �
�/�E�P�M$Qj;j �UR�M����P�E�P�Il�����M �U ��E�M��U�P�E�M�d�    Y��]�  ����������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P�����3�P�E�d�    �M�h�   h���EP�MQ�UR�EP� �����h�   h���M$Q蝯�����U�R�M�����E�E�E��E�    �M�Q�qc�����E��E������M���`���U�R�E$��Pjj �MQ�UR�E�P�������M �U ��E �8 uj �M�������Q�M���e���Ѓ�:t�E ����U �
�2�E�P�M$��Qj;j �UR�M諥��P�E�P谑�����M �U ��E �8 uj �M藐����Q�M��e���Ѓ�:t�E ����U �
�/�E�P�M$Qj;j �UR�M�G���P�E�P�L������M �U ��E�M��U�P�E�M�d�    Y��]�  ����������������������������������������������������������������������������������������������������������������������������U����M�hn  h���EP�MQ�UR�EP�h�����ho  h���M$Q茭�����U��BPj �MQ�UR��������E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U����M�hn  h���EP�MQ�UR�EP�/�����ho  h���M$Q�̬�����U��BPj �MQ�UR�>������E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U��j�h�d�    P�����3�P�E�d�    �M�h�  h���EP�MQ�UR�EP�ɩ����h�  h���M$Q�������U�R�M�e����E�E�E��E�    �M�Q�Y������E��E������M��]���E�    �U�R�E�Ph�  j �MQ�UR�E�P�-g�����M �U ��E ���u6�}�l  |�U���l  �U���}��   ~�E ����U �
�E$�M��H�U�E��M�J�E�M�d�    Y��]�  ��������������������������������������������������������������������������������U��j�h�d�    P�����3�P�E�d�    �M�h�  h���EP�MQ�UR�EP�Д����h�  h���M$Q�m������U�R�M�����E�E�E��E�    �M�Q�A^�����E��E������M��[���E�    �U�R�E�Ph�  j �MQ�UR�E�P��������M �U ��E ���u6�}�l  |�U���l  �U���}��   ~�E ����U �
�E$�M��H�U�E��M�J�E�M�d�    Y��]�  ��������������������������������������������������������������������������������U����M��E�    �E��HQ�M�k����U����U��E��]� ���������������U����M��E�    �E��HQ�M�+����U����U��E��]� ���������������U����M��E�    �E��HQ�M�����U����U��E��]� ���������������U����M��E�    �E��HQ�M諟���U����U��E��]� ���������������U��Q�M�j{hP��EP�MQ�_������U+U����R�EP�є������]� ���������������������U��Q�M�j{hP��EP�MQ��e�����U+U����R�EP联������]� ���������������������U����M�hq  h ��EP�MQ��z����hr  h ��UR�EP�u�����M�U��E �M��U�;Eu	�E�    ��E�   �M��M�U�;E��   �M �;U��   �E��P�MQ�U�E+P�M�R�E �Q�������E��U��U��}��t�}��t�}� t�4�E�M��E��]�   �V�U ����u�U�P�ͅ�������E��}��u�E�    �M�U��E��M ����E ��E�    �8����E��]� ����������������������������������������������������������������������������������U����M�h�  h ��EP�MQ�Ty����h�  h ��UR�EP��u�����M�U��E �M��U�;Eu	�E�    ��E�   �M��M�U�;E��   �M �;U��   �E��P�MQ�U�E+P�M�R�E �Q�Z������E��U��U��}��t�}��t�}� t�4�E�M��E��]�   �V�U ����u�U�P�=��������E��}��u�E�    �M�U��E��M ����E ��E�    �8����E��]� ����������������������������������������������������������������������������������U��Q�M�hk  h ��EP�MQ�~����hl  h ��UR�~������E���P�MQ�UR�EP��o������]� ������������������������U����M��E���P�MQ��q�������E#�t	�E�   ��E�    �E���]� �������������������������������U��Q�M�h�
  h ��EP�MQ�a����h�
  h ��UR讨�����E���P�MQ�UR�EP�"o������]� ������������������������U����M��E���P�MQ�q�������E#�t	�E�   ��E�    �E���]� �������������������������������U����M�h�  h ��EP�MQ�$v�����U��E��E�    �M�M��U�;U��   �E�;E��   �M��Q�U�R�E+E�P�M�Q�U�R�i������E��E��E�}��t�}��t�}� t�$�E��F�E��A�M���u�U�R�\��������E��}��u�E�    �E�E��E��M���M��a����E��]� ����������������������������������������������������������������U����M�h�  h ��EP�MQ�u�����U��E��E�    �M�M��U�;U��   �E�;E��   �M��Q�U�R�E+E�P�M�Q�U�R�I������E��E��E�}��t�}��t�}� t�$�E��F�E��A�M���u�U�R�<��������E��}��u�E�    �E�E��E��M���M��a����E��]� ����������������������������������������������������������������U��Q�M��   ��]�����������������U��Q�M��   ��]�����������������U��Q�M��EP�MQ�M��QU����]� �����������������U��Q�M�h�  h ��EP�MQ�Lz����h�  h ��UR�ِ������E���E�M���M�U;Ut�EP�M�R�M���T���M��ˋE��]� �����������������������������������������U��Q�M��EP�MQ�M��V����]� �����������������U��Q�M�h�
  h ��EP�MQ�/]����h�
  h ��UR�	�������E���E�M���M�U;Ut�EP�M�R�M��$V���M��ˋE��]� �����������������������������������������U��Q�M��E��H$�U�
�E��]� ���������������������U��Q�M��E��H$�U�
�E��]� ���������������������U����M��E�    �E��HQ�M�*[���U����U��E��]� ���������������U����M��E�    �E��HQ�M�u���U����U��E��]� ���������������U��Q�M������]� ����������������U��Q�M������]� ����������������U��� ���3ŉE��M�h�  h ��EP�MQ�w����h�  h ��UR�EP�p������M�U��E �M��U�;Eu	�E�    ��E�   �M�M�U�;E�  �M �;U�   �8����M �U+;�]�E��P�MQ�U��Q�U �P��������E��}� }�   �   �!�M����E��M �U��E ��E�    �   �M��U��E��P�MQ�U��Q�U�R蚟�����E��}� }	�   �]�S�E �M+;M�}�U�E���E��A�7�M�Q�U�R�E �Q�Z�����U����M��U �E��M ��E�    ������E�M�3���o����]� ����������������������������������������������������������������������������������������������������������U��� ���3ŉE��M�h�  h ��EP�MQ�SY����h�  h ��UR�EP�`������M�U��E �M��U�;Eu	�E�    ��E�   �M�M�U�;E�  �M �;U�   �(����M �U+;�]�E��P�MQ�U��Q�U �P�������E��}� }�   �   �!�M����E��M �U��E ��E�    �   �M��U��E��P�MQ�U��Q�U�R芝�����E��}� }	�   �]�S�E �M+;M�}�U�E���E��A�7�M�Q�U�R�E �Q�rX�����U����M��U �E��M ��E�    ������E�M�3��m����]� ����������������������������������������������������������������������������������������������������������U��Q�M��E��H �U�
�E��]� ���������������������U��Q�M��E��H �U�
�E��]� ���������������������U����M��E�    �E��HQ�M��U���U����U��E��]� ���������������U����M��E�    �E��HQ�M�vp���U����U��E��]� ���������������U��j�h0d�    P��d���3ŉE�P�E�d�    �M��E�P�M��p���E��M��M��E�    �U�R��|�����E��E������M��I���E�P�   k��¨�R�   k� ����Q�M��Ë���E� �E�    �M �p{���Ѕ�u+j �M ��\��� �   k�
�L�;�u�E��U����U��M �~����E��E��E��	�M����M��U�;U�s&�E�P�M �s\��f���R�E�P�h�������
s�ɋM�+M�Q�U�R�M �F\��P�M�趒���E�   �M���z������t�   k� �D�Pj�M�赗���   k� �D�P���̉e��U�R�w���E��E�P�MQ�UR�EP�MQ�UR�EP�M��)b���E������M���Z���E�M�d�    Y�M�3��j����]� ����������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��t���3ŉE�P�E�d�    �M��E� ���] ����Au�E��E ���] �E�    �	�E���
�E��E ������u�}��  s�E �5���] �Ѓ��E �$h�j(�M�Q�ք�����E��}� }�U�E��M�J�E��   �U�R�M�
n���E��E��E��E�    �M�Q��y�����E��E������M��F��j0�M���Y��f�E�j �U�R�M��F���E�   j �M��]��P�E��L�Q�   k� �L�Q�M�貈���U�R�E�P�M��l����M�Q���̉e��U�R�Nu���E��E�P�MQ�UR�EP�MQ�UR�EP�M���_���E������M��X���E�M�d�    Y�M�3��Uh����]�  ������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��d���3ŉE�P�E�d�    �M��E�P�M�jl���E��M��M��E�    �U�R��G�����E��E������M��E���E�P�   k����R�   k� ���Q�M��Y���E� �E�    �M �K���Ѕ�u+j �M �%I��� �   k�
�L�;�u�E��U����U��M �5����E��E��E��	�M����M��U�;U�s&�E�P�M ��H��f���R�E�P��������
s�ɋM�+M�Q�U�R�M �H��P�M��o^���E�   �M���J������t�   k� �D�Pj�M������   k� �D�P���̉e��U�R�3R���E��E�P�MQ�UR�EP�MQ�UR�EP�M�趋���E������M���r���E�M�d�    Y�M�3��f����]� ����������������������������������������������������������������������������������������������������������������������������������U��j�h d�    P��t���3ŉE�P�E�d�    �M��E� ���] ����Au�E��E ���] �E�    �	�E���
�E��E ������u�}��  s�E �5���] �Ѓ��E �$h�j(�M�Q�F������E��}� }�U�E��M�J�E��   �U�R�M�zi���E��E��E��E�    �M�Q��D�����E��E������M��-B��j0�M��`���f�E�j �U�R�M������E�   j �M��~n��P�E��L�Q�   k� �L�Q�M�� V���U�R�E�P�M�襕���M�Q���̉e��U�R��O���E��E�P�MQ�UR�EP�MQ�UR�EP�M��v����E������M��p���E�M�d�    Y�M�3���c����]�  ������������������������������������������������������������������������������������������������������������������U���P���3ŉE��M��EP�M�v���Phؗ�M�Q�U�R�x`����Pj@�E�P�n~����P�M�Q�UR�EP�MQ�UR�EP�M�Q�R���� �E�M�3���b����]� �����������������������������������U���P���3ŉE��M��EP�M�ֈ��Phܗ�M�Q�U�R��_����Pj@�E�P��}����P�M�Q�UR�EP�MQ�UR�EP�M�Q��Q���� �E�M�3��6b����]� �����������������������������������U���   ���3ŉE���`����M�$�����T�����X�����X��� 0|	��T��� w%�M����%    uǅh���   ǅl���    ��M�׈����h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M�X���% 0  =    �  �E�@v�E������D��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E������u��x����  s�E�5���]���E��s����Aud���t�����
��t����}� |M	��|���
rB�Й�]����u2��t����  s&�E����]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M����Pj �E�P��`���Q�&e����Pjl�U�R�{����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P�����,�E�M�3��e_����]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE���`����M�ą����T�����X�����X��� 0|	��T��� w%�M謄��%    uǅh���   ǅl���    ��M�w�����h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M�����% 0  =    ��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E������u��x����  s�E�5���]���E��s����Aud���t�����
��t����}� |M	��|���
rB�Й�]����u2��t����  s&�E����]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M�ւ��PjL�E�P��`���Q��a����Pjl�U�R��w����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P�m|����,�E�M�3��\����]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���H���3ŉE��M��EPh�j@�M�Q�v����P�U�R�EP�MQ�UR�EP�MQ�U�R�J���� �E�M�3��[����]� �����������������������������U���P���3ŉE��M��E P�MQ�M����Ph���U�R�E�P�X����Pj@�M�Q�
v����P�U�R�EP�MQ�UR�EP�MQ�U�R�J���� �E�M�3��rZ����]� �����������������������������������������������U���P���3ŉE��M��E P�MQ�M�b���Ph��U�R�E�P�dW����Pj@�M�Q�Zu����P�U�R�EP�MQ�UR�EP�MQ�U�R�oI���� �E�M�3���Y����]� �����������������������������������������������U��j�hsd�    P��   ���3ŉE�VP�E�d�    �M�h�  hx��EP�F�����M���% @  u4�MQ�UR�EP�MQ�UR�EP�M���M��B$�ЋE��  ��  ��p���Q�M�]���E��U���|����E�    ��|���P��c�����E��E�������p����d6���M�蜇���E�   �M��t%�U�R�M��>���E��E�P�M���o���M���H���#�M�Q�M���P���E��U�R�M��o���M��H���M��c����t�����x�����x��� |:	��t��� v/�M�c�����M�����;�v�M�c�����M������+��u���E�    �E��E��M�<~��%�  ��@t6�M�Q�UR�EP�MQ��`���R�E�P�<�������P�M�U�E�    �M�虃��P�M��\��P�EP�MQ��h���R�E�P��b������P�M�Uj j �M��H���E�P�MQ�UR�EP�MQ�U�R�ń�����E������M��G���E�M�d�    Y^�M�3��'W����]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������U���P���3ŉE��M��EP�M�|��Phؗ�M�Q�U�R��k����Pj@�E�P�q����P�M�Q�UR�EP�MQ�UR�EP�M�Q�u���� �E�M�3��V����]� �����������������������������������U���P���3ŉE��M��EP�M�|��Phܗ�M�Q�U�R�Yk����Pj@�E�P��p����P�M�Q�UR�EP�MQ�UR�EP�M�Q�u���� �E�M�3��fU����]� �����������������������������������U���   ���3ŉE���`����M�T|����T�����X�����X��� 0|	��T��� w%�M�<{��%    uǅh���   ǅl���    ��M�|����h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M�z��% 0  =    �  �E�@v�E������D��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E������u��x����  s�E�5���]���E��s����Aud���t�����
��t����}� |M	��|���
rB�Й�]����u2��t����  s&�E����]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M�My��Pj �E�P��`���Q�nJ����Pjl�U�R�En����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P�g����,�E�M�3��R����]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE���`����M��x����T�����X�����X��� 0|	��T��� w%�M��w��%    uǅh���   ǅl���    ��M�x����h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M�(w��% 0  =    ��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E������u��x����  s�E�5���]���E��s����Aud���t�����
��t����}� |M	��|���
rB�Й�]����u2��t����  s&�E����]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M�v��PjL�E�P��`���Q�'G����Pjl�U�R��j����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P��c����,�E�M�3��NO����]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���H���3ŉE��M��EPh�j@�M�Q��i����P�U�R�EP�MQ�UR�EP�MQ�U�R��m���� �E�M�3��@N����]� �����������������������������U���P���3ŉE��M��E P�MQ�M�Bt��Ph���U�R�E�P�c����Pj@�M�Q�:i����P�U�R�EP�MQ�UR�EP�MQ�U�R�Bm���� �E�M�3��M����]� �����������������������������������������������U���P���3ŉE��M��E P�MQ�M�s��Ph��U�R�E�P��b����Pj@�M�Q�h����P�U�R�EP�MQ�UR�EP�MQ�U�R�l���� �E�M�3���L����]� �����������������������������������������������U��j�h�d�    P��   ���3ŉE�VP�E�d�    �M�h�  hx��EP�)v�����M�r��% @  u4�MQ�UR�EP�MQ�UR�EP�M���M��B$�ЋE��  ��  ��p���Q�M��P���E��U���|����E�    ��|���P�3*�����E��E�������p����)���M���Z���E�   �M��t%�U�R�M��~v���E��E�P�M��s^���M��vX���#�M�Q�M���5���E��U�R�M��N^���M��QX���M�W����t�����x�����x��� |:	��t��� v/�M��V�����M��q��;�v�M��V�����M��tq��+��u���E�    �E��E��M�lq��%�  ��@t6�M�Q�UR�EP�MQ��`���R�E�P��h������P�M�U�E�    �M��q��P�M��"`��P�EP�MQ��h���R�E�P�T������P�M�Uj j �M�<���E�P�MQ�UR�EP�MQ�U�R�Kh�����E������M��1W���E�M�d�    Y^�M�3��WJ����]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hd�    P��T���3ŉE�P�E�d�    �M�h&  h���EP�6����h'  h���MQ��W�������U���E�f��f�M�M��<X���E�    �U$��uf�E �   ��f�D��#f�U$�   ��f�T�f�M �   k�f�L��E�   ��M���M�j �U�R�M��Gz���M����LG��P�EP�M�Q�M���n��P�U�R�M��3j���E��E��E��E��M���3��P��b�����E��}� v	�E�   ��E�    �M��M��E� �M���6���Uǅ�t��i����EP�MQ�U�R�M��\R��Pj�M��QR��P�EP��]�����E������M���T���E�M�d�    Y�M�3���G����]�  �����������������������������������������������������������������������������������������������������������������������U��j�h`d�    P��T���3ŉE�P�E�d�    �M�h�  h���EP��p����h�  h���MQ�U�������U���E�f��f�M�M��V���E�    �U$��uf�E �   ��f�D��#f�U$�   ��f�T�f�M �   k�f�L��E�   ��M���M�j �U�R�M��x���M����E��P�EP�M�Q�M��l��P�U�R�M��h���E��E��E��E��M��1��P�`�����E��}� v	�E�   ��E�    �M��M��E� �M��4���Uǅ�t��i����EP�MQ�U�R�M��,P��Pj�M��!P��P�EP�8�����E������M��R���E�M�d�    Y�M�3���E����]�  �����������������������������������������������������������������������������������������������������������������������U��Q�M�ht  h ��EP�MQ�K�����	�U���U�E;Et�M�R�EP�M��k���ȅ�u�ҋE��]� ����������������������U��Q�M�h�
  h ��EP�MQ��.�����	�U���U�E;Et�M�R�EP�M���?���ȅ�u�ҋE��]� ����������������������U��Q�M�h}  h ��EP�MQ�J�����	�U���U�E;Et�M�R�EP�M���j���ȅ�t�ҋE��]� ����������������������U��Q�M�h�
  h ��EP�MQ��-�����	�U���U�E;Et�M�R�EP�M��
?���ȅ�t�ҋE��]� ����������������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M��E���P�MQ�]������]� ���������������U��Q�M�h�  h ��EP�MQ�,I�����	�U���U�E;Et�M���Q�U�P�]]�����Mf��ыE��]� �������������������������������������U��Q�M�h�
  h ��EP�MQ�_,�����	�U���U�E;Et�M���Q�U�P��\�����Mf��ыE��]� �������������������������������������U��Q�M��E���P�MQ�\������]� ���������������U��Q�M��E���P�MQ�Rp������]� ���������������U��Q�M�h�  h ��EP�MQ��G�����	�U���U�E;Et�M���Q�U�P��o�����Mf��ыE��]� �������������������������������������U��Q�M�h�
  h ��EP�MQ��*�����	�U���U�E;Et�M���Q�U�P�so�����Mf��ыE��]� �������������������������������������U��Q�M��E���P�MQ�"o������]� ���������������U��j�h�d�    P��\���3ŉE�VP�E�d�    �M��E�    jhhP��EP�MQ�sF�����M���n���E�    �U+U���Ũ}� ��   �E�P�M��_���M���Q�UR�EP�M�Q�M��1���E��U��U��E��M��C�����M��k���FP�M�Q�M��1���E��U��U��E��M���B��P�(&�����E̍M��Mk��9E�w	�E�   ��E�    �EȈE��E��M��:%���E� �M��.%���MӅ�t��5����U�R�M���^���E�P�M�A���Mă��M��E������M��?/���E�M�d�    Y^�M�3���>����]� ��������������������������������������������������������������������������������������������������U��j�hd�    P��\���3ŉE�VP�E�d�    �M��E�    jhhP��EP�MQ�F(�����M��%M���E�    �U+U���Ũ}� ��   �E�P�M��`���M���Q�UR�EP�M�Q�M��f_���E��U��U��E��M�� )�����M���c���FP�M�Q�M��7_���E��U��U��E��M���(��P�Wj�����E̍M��c��9E�w	�E�   ��E�    �EȈE��E��M���+���E� �M��+���MӅ�t��5����U�R�M��G_���E�P�M��T���Mă��M��E������M���I���E�M�d�    Y^�M�3���<����]� ��������������������������������������������������������������������������������������������������U����M��E�    �E��HQ�M�%���U����U��E��]� ���������������U����M��E�    �E��HQ�M�@���U����U��E��]� ���������������U������3ŉE��M�h�  h ��EP�MQ�*Y�����U�E��E�    �M��U�E��P�MQj �U�R�k�����E��}� 	�E�   �P�E����E��M�U+;U�}�E�M��E�   �)�}� ~#�U�R�E�P�M�R��%�����E�M��U�
�E�M�3��A;����]� ��������������������������������������������������������������U������3ŉE��M�h�  h ��EP�MQ�X�����U�E��E�    �M��U�E��P�MQj �U�R��i�����E��}� 	�E�   �P�E����E��M�U+;U�}�E�M��E�   �)�}� ~#�U�R�E�P�M�R��$�����E�M��U�
�E�M�3��1:����]� ��������������������������������������������������������������U��Q�M��EP�M��G5����]� ������U��Q�M�h�  h ��EP�MQ�F9����h�  h ��UR�5H������E���E�M���M�U;Ut�E�Q�M���4���Uf��ϋE��]� �����������������������������U��Q�M�h�
  h ��EP�MQ�8����h�
  h ��UR�?������E���E�M���M�U;Ut�E�Q�M���P���Uf��ϋE��]� �����������������������������U��Q�M��EP�M��P����]� ������U����M��E��x u	�E�   ��E�    �E���]������������������������U����M��E��x u	�E�   ��E�    �E���]������������������������U��Q�M��E�P�M��L,���M��Q�PP�M�]���E��]� ������������������U��Q�M��E�P�M��H���M��Q�PP�M�FX���E��]� ������������������U����  ]�������U����  ]�������U��Q�E��U�;�u	�E�   ��E�    �E���]����������������������U��Q�E��U�;�u	�E�   ��E�    �E���]����������������������U����M��E��H��u�M�����U�B��u�M����M��9 u�U�: t�E��8 t�M�9 u	�E�    ��E�   �E���]� ����������������������������������������U����M��E��H��u�M��^Z���U�B��u�M�KZ���M��9 u�U�: t�E��8 t�M�9 u	�E�    ��E�   �E���]� ����������������������������������������U��Q�M��E��H;Ms�M��/���UR�M��=���E���]� �����������������U����M��E��H;Ms�M���.���U��B+E;Ew�MQ�M��m=���L�} vF�M��)���U�P�E��M��Q+U�U�E�+EP�M�U��JP�M�Q�/<�����U�R�M��=���E���]� �����������������������������������U��Q�M��E��H;Ms�M��L���UR�M��'���E���]� �����������������U����M��E��H;Ms�M��nL���U��B+E;Ew�MQ�M��L'���L�} vF�M��UE���U�P�E��M��Q+U�U�E�+EP�M�U��JP�M�Q�B�����U�R�M���&���E���]� �����������������������������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��E���M��B$�Ћ�]���������U��Q�M��E���M��B$�Ћ�]���������U����M��E�P�M����P�M�a���E��]� ���������U����M��E�P�M����P�M�CL���E��]� ���������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P �ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P �ҋE��]�  �������������������U��Q�M��E��H���]��������������U��Q�M��E��H���]��������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E��H;Ms�M���(���U��P�+B;Ew�M��M���} vx�M��QU�U�j �E�P�M��Y���ȅ�tW�U��B+EP�M��#���M�HR�M��#���M�H�E�BQ�66�����UR�EP�MQ�M��5���U�R�M��7���E���]� �����������������������������������������������������U����M��E��H;Ms�M��F���U����+B;Ew�M��]���} vx�M��QU�U�j �E�P�M��\"���ȅ�tW�U��B+EP�M��N?���M�HR�M��??���M�H�E�BQ�I�����UR�EP�MQ�M�����U�R�M��� ���E���]� �����������������������������������������������������U��Q�M��EP�MQ�U���M��P�ҋ�]� ������������U��Q�M��EP�MQ�U���M��P�ҋ�]� ������������U��Q�E���u	�E�    ��UR�.8�����E��E���]��������������������U��Q�E���u	�E�    ��UR��7�����E��E���]��������������������U��Q�M��E�P��-������]����������U��Q�M��E�P�������]����������U��Q�M�������]�����������������U��Q�M�������]�����������������U��M�;��]����U��M�P��]����U����M��E�P�M����������E��}�w	�E�   �	�M����M�E��]�������������������U����M��E�P�M�������D���E��}�w	�E�   �	�M����M�E��]�������������������U��Q�} u�E�E���MQ�UR�EP�S�����E��E���]�����������������U��Q�} u�E�E���MQ�UR�EP�wS�����E��E���]�����������������U��j�hYd�    P��X���3ŉE�P�E�d�    �M��E�    �E��8 u)�M��
W���E��M��M��E�    �U����U��E��E��(�M��	���\;��P�M��1N���E��U����U��E��E��M��M��U�R�M�`���E����E��M���t�e���M�����E������U���t�e���M�����E�M�d�    Y�M�3��@*����]� �������������������������������������������������������������U��Q�M��EP�MQ�U���M��P8�ҋ�]� ������������U��Q�M��EP�MQ�U���M��P8�ҋ�]� ������������U��Q�M��EP�M���M��B,�ЋE��]� ���������������U��Q�M��EP�M���M��B,�ЋE��]� ���������������U����M��E�    �EP�M���M��B �ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B �ЋM����M��E��]� �������������U��Q�M��EP�M���M��B(�ЋE��]� ���������������U��Q�M��EP�M���M��B(�ЋE��]� ���������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E��H;Mr�M�S��;Es�M��!���U��B+E;Es�M��Q+U�U�M�S��+E�E��E�;Es�M��M���+U�E��H+M;�w�M��E���U��B+E+E�E��M��QU+U�U�E��H;M�sj �U�R�M��kQ���E�;Ete�M�Q�M��j���U�P�M�HR�M��U���M�H�E�BQ�.�����UR�M�����M�HR�M��%���M�HR�G������  �E;Ewe�MQ�M������U�PP�M������M�HR�-�����E�P�M������M�H�E�BQ�M�����U�P�M�HR�q-�����|  �E;Ewe�M�Q�M�����U�P�M�HR�M��{���M�H�E�BQ�.-�����UR�M��Z���M�HR�M��K���M�HR�-�����  �EE;Ewk�M�Q�M�� ���U�P�M�HR�M�����M�H�E�BQ�,�����UR�M������MM+M�HR�M������M�HR�,�����   �EP�M�����M�HR�M�����M�HR�_,�����E�P�M�����M�H�E�BQ�M��v���U�P�M�HR�),�����E+EP�M��R���M�H�E�BQ�M��=���U�P�M�HR��+�����E�P�M���,���E���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��} th�  h ��EP��+�����MQ�M��K���Ѕ�t-�EP�M������M+���Q�U�R�EP�MQ�M��G���5  �U��B;Es�M������M��Q+U;Us�E��H+M�M���+U�E��H+M;�w�M��hA���U��B+E+E�E��M;Ms6�U�R�M��o���M�H�E�BQ�M��Z���U�P�M�HR�*�����} w
�} ��   �E��HM+M�M�j �U�R�M��M������ti�M;Ms6�U�R�M������M�H�E�BQ�M������U�P�M�HR�)�����EP�MQ�M������U�PP�������M�Q�M��l*���E���]� ����������������������������������������������������������������������������������������������������������������U��j�h�d�    P��   ���3�P�E�d�    �M��E�   �E,P�M �(���ȅ���   ���̉e��UR�O���EȋEȉE��E����̉e��UR�nO���E��E��%(�����EЋE�P��p���Q�M��D���E��U��U��E����̉e��E�P�+O���E؋M؉M��E����̉e��UR�O���E��E���'�����E�E�P�M������E���p���������   �M Q�M,��!��P�M �$��P���̉�|����UR�N���E�E�E��E����̉e��UR�N���E��E��J'�����E�E�P��d���Q�M��i���E܋U܉U��E����̉e��E�P�PN���E̋M̉M��E�	���̉e��UR�2N���E��E���&�����EċE�P�M��/���E���d��������M��M��E��M�6���E��M�*���E� �M �����E������M,�����E��M�d�    Y��]�0 ��������������������������������������������������������������������������������������������������������������������������������������������������U����M��E��H;Mr�M�5E��;Es�M���6���U��B+E;Es�M��Q+U�U�M�E��+E�E��E�;Es�M��M���+U�E��H+M;�w�M��)M���U��B+E+E�E��M��QU+U�U�E��H;M�sj �U�R�M��_���E�;Ete�M�Q�M��V/���U�P�M�HR�M��A/���M�H�E�BQ�K	�����UR�M�.���M�HR�M��/���M�HR�m������  �E;Ewe�MQ�M���.���U�PP�M���.���M�HR�������E�P�M��.���M�H�E�BQ�M��.���U�P�M�HR������|  �E;Ewe�M�Q�M��|.���U�P�M�HR�M��g.���M�H�E�BQ�q�����UR�M��F.���M�HR�M��7.���M�HR�G�����  �EE;Ewk�M�Q�M��.���U�P�M�HR�M���-���M�H�E�BQ������UR�M���-���MM+M�HR�M���-���M�HR�������   �EP�M��-���M�HR�M��-���M�HR������E�P�M��w-���M�H�E�BQ�M��b-���U�P�M�HR�l�����E+EP�M��>-���M�H�E�BQ�M��)-���U�P�M�HR�3�����E�P�M������E���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��} th�  h ��EP�e �����MQ�M��@���Ѕ�t-�EP�M���+���M+���Q�U�R�EP�MQ�M��<G���5  �U��B;Es�M��2���M��Q+U;Us�E��H+M�M���+U�E��H+M;�w�M��I���U��B+E+E�E��M;Ms6�U�R�M��[+���M�H�E�BQ�M��F+���U�P�M�HR�P�����} w
�} ��   �E��HM+M�M�j �U�R�M���������ti�M;Ms6�U�R�M���*���M�H�E�BQ�M���*���U�P�M�HR�������EP�MQ�M��*���U�PP�������M�Q�M��{���E���]� ����������������������������������������������������������������������������������������������������������������U��j�h�d�    P��   ���3�P�E�d�    �M��E�   �E,P�M �D���ȅ���   ���̉e��UR������EȋEȉE��E����̉e��UR�����E��E���	�����EЋE�P��p���Q�M��:���E��U��U��E����̉e��E�P�{����E؋M؉M��E����̉e��UR�]����E��E��	�����E�E�P�M��w����E���p��������   �M Q�M,�3��P�M �:��P���̉�|����UR�����E�E�E��E����̉e��UR������E��E��"	�����E�E�P��d���Q�M��39���E܋U܉U��E����̉e��E�P�����E̋M̉M��E�	���̉e��UR�����E��E��������EċE�P�M�����E���d�������M��M��E��M������E��M������E� �M �~���E������M,�o���E��M�d�    Y��]�0 ��������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M�j �EP�M�������]� ���������������������U��Q�M��E��M;Hw�UR�M��%����EP�M��U+QR�M��B����]� �������������������U��Q�M�j �EP�M��3����]� ���������������������U��Q�M��E��M;Hw�UR�M��t����EP�M��U+QR�M���F����]� �������������������U����M��M��v"���E��U�}� |�}� v�M��a���P�q����f�E���E���M��B��f�E�f�E���]����������������������������U����M��M��f?���E��U�}� |�}� v�M��{;��P�h����f�E���E���M��B��f�E�f�E���]����������������������������U����M��E�P�M�Q�#?����P�M�����E��]� ���������������������U����M��E�P�M�Q�D����P�M�G3���E��]� ���������������������U��Q�M��E�P�M�B���E��]� ��������������������U��Q�M��E�P�M�-���E��]� ��������������������U��EP�M�U����E]�������������U��EP�M�W>���E]�������������U����M��M��v ���E��U�}� |�}� v�M����P�q����f�E���E���M��B��f�E�f�E���]����������������������������U����M��M��f=���E��U�}� |�}� v�M��>��P�h
����f�E���E���M��B��f�E�f�E���]����������������������������U��Q�M��E��@��]����������������U��Q�M��E��@��]����������������U����M��M��=���E�U��}� |/�}� v'�M�������E�E�f�Mf��U�R�A����f�E��!�EP�/������Q�U���M��P��f�E�f�E���]� �����������������������������������������U����M��M�����E�U��}� |/�}� v'�M������E�E�f�Mf��U�R�	����f�E��!�EP��������Q�U���M��P��f�E�f�E���]� �����������������������������������������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Ef� ]������U��Ef� ]������U��Ef� ]������U��Ef� ]������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��EP�M���M��B0�Ћ�]� �����������������U��Q�M��EP�MQ�UR�E���M��B,�Ћ�]� ����������U��Q�M��EP�MQ�UR�E���M��B,�Ћ�]� ����������U��Q�M��EP�M���M��B0�Ћ�]� �����������������U��E��P�MQ�UR�f�����]����������������������U��E��P�MQ�UR������]����������������������U��Q�E�E���M����M��U���U�} v�E�f�Mf��܋E��]��������������������������U��Q�EP�MQ������E��U�R�EP�MQ�UR�EP�MQ�e�����E��]������������������U��Q�EP�M�Q�������UR�E�P������M�Q�U�R�EP�MQ�UR�EP�MQ��������E��]��������������������������������U����M������E���E�M;Mt�U�P�M�6�����=���ϋM�U��E�A�E]������������������������U��EP�MQ�UR�EP�MQ�P
�����E]�������������U����M��E��H(��t�U�B�E��	�M�Q�U��E���,Pj �M�Q��������U��B�E�H.��v	�E��a�	�U�B �E�M���,Qj �U�R�������M��A�U�B/��v	�E��	�M�Q$�U��E���,Pj �M�Q�r������U��B�E���,Pj �   k� �E�H�R�������M��A�U���,Rj �   k� �U�B�Q�������U��B��]� ���������������������������������������������������������������������������������U���4���3ŉE�VW�M̍E�P�M����}̃��   ���M̃�Qj �M�4���P�w������ỦB�Ẽ�Pj �M�D���P�W������M̉A�Ũ�Rj hX��;������M̉A_^�M�3������]� ��������������������������������������������������U��Q3��E��E���]�����������������U��E]���������U��EP�MQ�UR�EP�MQ�L0����]����������������U��EP�MQ�UR�EP�MQ��5����]����������������U��Q�E���]������U��E]���������U��j�hd�    P��`���3�P�E�d�    �M��E�   ���̉eȍEP�H���E�M�M��E����̉e��UR�*���E�E�E��E��M�Q�M��J����E�U�U��E����̉e��E�P�0���E܋M܉M��E��U�R�M��!���E؋E؉E��E����̉e��U�R�����E��E��M���$���EЋEЉE��E��M��D���E��M��8���E� �M�,���E������M����E̋M�d�    Y��]� �������������������������������������������������������������������������������������U��Q�E;Eu�M�U��E�A�E�{�yhQ  h ��MQ�UR�%����hR  h ��EP�������MQ�UR�>�����E��E�P�MQ�UR�EP�O	����P�MQ�B	����P�UR�X	�����E��]���������������������������������������������������U��j�hHd�    P��$���3�P�E�d�    j �M��)����E�    �p��E�P��A����E�M�Q�M�y���E�}� t�n�}� t�U��U��`�EP�M�Q�\ �������uhDq�M��>���hPP�U�R�d���.�E��E�M��p��U��U�E��M�B�ЋM�Q�&�����U�U��E������M�����E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hxd�    P��$���3�P�E�d�    j �M�������E�    �t��E�T������E�M�Q�M�9���E�}� t�n�}� t�U��U��`�EP�M�Q���������uhDq�M������hPP�U�R�$���.�E��E�M��t��U��U�E��M�B�ЋM�Q��$�����U�U��E������M��v���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M������E�    �x��E�X�������E�M�Q�M�����E�}� t�n�}� t�U��U��`�EP�M�Q���������uhDq�M�����hPP�U�R�����.�E��E�M��x��U��U�E��M�B�ЋM�Q�#�����U�U��E������M��6���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M��i����E�    �|��E�\������E�M�Q�M����E�}� t�n�}� t�U��U��`�EP�M�Q��$�������uhDq�M��~���hPP�U�R����.�E��E�M��|��U��U�E��M�B�ЋM�Q�D"�����U�U��E������M������E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hd�    P��$���3�P�E�d�    j �M��)����E�    ����E�d��A����E�M�Q�M�y���E�}� t�n�}� t�U��U��`�EP�M�Q��������uhDq�M��>���hPP�U�R�d���.�E��E�M�����U��U�E��M�B�ЋM�Q�!�����U�U��E������M�����E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h8d�    P��$���3�P�E�d�    j �M�������E�    ����E�`������E�M�Q�M�9���E�}� t�n�}� t�U��U��`�EP�M�Q��$�������uhDq�M������hPP�U�R�$���.�E��E�M�����U��U�E��M�B�ЋM�Q�������U�U��E������M��v���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hhd�    P��$���3�P�E�d�    j �M������E�    ����E�h�������E�M�Q�M�����E�}� t�n�}� t�U��U��`�EP�M�Q�V��������uhDq�M�����hPP�U�R�����.�E��E�M�����U��U�E��M�B�ЋM�Q������U�U��E������M��6���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M��i����E�    ����E�l������E�M�Q�M����E�}� t�n�}� t�U��U��`�EP�M�Q��������uhDq�M��~���hPP�U�R����.�E��E�M�����U��U�E��M�B�ЋM�Q�D�����U�U��E������M������E܋M�d�    Y��]��������������������������������������������������������������������������U��Q�M��EP�M�����E���]� ��������������������U��j�h�d�    PQ���3�P�E�d�    �M��EP�M�����E�    �M��d��U��E�B(�MQ�UR�M��n����E������E��M�d�    Y��]� �����������������������������������������U��Q�M��EP�M�������M��U�B�A�E���]� ������������������������U��Q�M��M�����E��@    �E���]�����������������U��Q�M��EP�M��"���E���]� ��������������������U��j�h�d�    P�����3�P�E�d�    �M�M��"��P�M��S����E�    j j �M������EP�MQ�M��^���E������E�M�d�    Y��]� �����������������������������������������U��j�h(	d�    PQ���3�P�E�d�    �M��EP�M�������E�    �M�����UR�M��,���E������E��M�d�    Y��]� ���������������������������������������U��j�hX	d�    PQ���3�P�E�d�    �M��EP�M�� !���E�    �M����UR�M���*���E������E��M�d�    Y��]� ���������������������������������������U��j�h�	d�    PQ���3�P�E�d�    �M��EP�M������E�    �M��,��UR�M������E������E��M�d�    Y��]� ���������������������������������������U��j�h�	d�    PQ���3�P�E�d�    �M��EP�M������E�    �M��H��UR�M�������E������E��M�d�    Y��]� ���������������������������������������U��Q�M��EPj�MQ�UR�M�������E�� ��E���]� ����������������U��Q�M��EPj �MQ�UR�M������E�� ���E���]� ����������������U��j�h�	d�    PQ���3�P�E�d�    �M��EP�M������E�    �M��$��UR�M��;����E������E��M�d�    Y��]� ���������������������������������������U��j�h#
d�    PQ���3�P�E�d�    �M��EP�M��u����E�    �M��X�j �M����l���E��UR�M��5����E������E��M�d�    Y��]� ��������������������������������������U��Q�M��E�� d��M��X"���M�������]�������������U��Q�M��E�� ���M��QR�������M��F�����]����������������������U��Q�M��E�� ��M������]���������������������U��Q�M��E�� ,��M��������]���������������������U��Q�M��E�� H��M�������]���������������������U��Q�M��E�� ��M��	����]���������������������U��Q�M��E�� ���M�������]���������������������U��Q�M��E�� $��M��8'���M������]�������������U��Q�M��E�� X��M�������M��������]����������U��Q�M��EP�M������E���]� ��������������������U��Q�M��EP�M�������M��U�B�A�E���]� ������������������������U����M��E�;E��   j j�M������3�t�U�R�M���P�M��d���E�P�M���P�M�Q�M����P�Z������Ѕ�t,���ĉe�P�M��������̉e�Q�M�����M��s�����UR������P�M��>����E���]� ���������������������������������������������������U����M��EP�M������M��U�A;Bu	�E�   ��E�    �E���]� ��������������������U����M��EP�M��"���ȅ�u	�E�   ��E�    �E���]� ���������������������������U��QV�M��M��g�����t-�E��x t$�M��R������k������M��A���p�M�;qw_jmh �h����������i��t3�u#hjhpjj jnh �j���������u�j jnh �h��h�k������U��B���M��A�E�^��]����������������������������������������������������������U��Q�M��E���]� ����������������U��Q�M��EP�M������M��U�A+B��]� �����������U��j�hX
d�    P�����3�P�E�d�    �M��E�    �E�P�M������E�    �MQ�M��}��P�M������U����U��E������M������E�M�d�    Y��]� ���������������������������������������������U��j�h�
d�    P�����3�P�E�d�    �M��EP�M�Q�M�����E�U�U��E�    �M������E��E������M�������E�M�d�    Y��]� ������������������������������������������U��j�h�
d�    P�����3�P�E�d�    �M��E�    �E�P�M������E�    �MQ�M�����P�M�����U����U��E������M��5����E�M�d�    Y��]� ���������������������������������������������U��QV�M��M��'�����tN�E��x tE�M��qu�M��	������"���;�r)�M���������������M������p�U��BE;�shh�   h �h��~�������i��t3�u&hjhpjj h�   h �j�m�������u�j h�   h �h��h�k������M��QU�E��P�E�^��]� �������������������������������������������������������������U��Q�M��EP�M�����E���]� ��������������������U��Q�M��E��P�M��&
����]� ���������������������U��Q�M��M������E��t�M�Q��������E���]� ��������������������U��Q�M��M������E��t�M�Q�������E���]� ��������������������U��Q�M��M��	����E��t�M�Q�O������E���]� ��������������������U��Q�M��M�������E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q��������E���]� ��������������������U��Q�M��M��d���E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q�O������E���]� ��������������������U��Q�M��M��	���E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q��������E���]� ��������������������U��QV�M��M��g�����t�M��[������M�Q���;�thh�   h �hh����������m��t3�u&h(nhpjj h�   h �j���������u�j h�   h �hx�h�o�����^��]� ���������������������������������������U��j�h-d�    P��x���3ŉE�P�E�d�    �E�    �} ��   �E�8 ��   ����E�jCh ��M�Qj�������E��E�    �}� tbj �U�R�M�R����E��E��E��E��MЃ��MЋM������P��|���������E��U��U��E�   �EЃ��EЋM�Q�M�����E���E�    �UȉU��E�   �E�M���E�   �UЃ�t�e����|�������E������EЃ�t�e���M��m����   �M�d�    Y�M�3�������]������������������������������������������������������������������������������������������U��j�h�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�jMh���M�Qj�p������E��E�    �}� t:j �M����P�M��|����E��U��U��E��E����E��M�Q�M��W����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]�����������������������������������������������������������������������������U��j�hd�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h�  h��M�Qj�-������E��E�    �}� t:j �M� ��P�M��9����E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��e���   �M�d�    Y��]��������������������������������������������������������������������������U��j�htd�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �m����E�h�  h��M�Qj��������E��E�    �}� t:j �M�Y���P�M�������E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��%���   �M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �-����E�h(  h��M�QjX�������E��E�    �}� t<jj �M����P�M������E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]������������������������������������������������������������������������U��j�hTd�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�h(  h��M�QjX�m������E��E�    �}� t<jj �M�����P�M��w����E��U��U��E��E����E��M�Q�M�����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]������������������������������������������������������������������������U��j�h�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h�   h|��M�QjD�-������E��E�    �}� t:j �M����P�M��9����E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��e���   �M�d�    Y��]��������������������������������������������������������������������������U��j�h4d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �m����E�h�  h|��M�Qj��������E��E�    �}� t:j �M�Y���P�M�������E��U��U��E��E����E��M�Q�M��Y���E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��%���   �M�d�    Y��]��������������������������������������������������������������������������U��j�hxd�    P�����3�P�E�d�    �M��E�P�M�����E�M�M��E�    �U�R�������E��E������M��@����	�E(���E(�M(�����   �E(���%uO�U(���U(j �E(�Q�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M���M��B$�Ћ�P�M�U�   �E(��� uB��M�q����UR�EP�]������ȅ�t�M�������RjH�M����������t���<j �M������Q�M��X����ЋE(�;�t�U ����M ����M����������UR�EP�������ȅ�t�U ����M ��U�E��M�J�E�M�d�    Y��]�$ �����������������������������������������������������������������������������������������������������������������������U���@���3ŉE��E܉EԋMQ�UR�����������t�[j �M������Q�M �+����E��Uۃ�+u�E�� +�Mԃ��MԋM������ �Uۃ�-u�E�� -�Mԃ��MԋM�����E� �UR�EP�������ȅ�t,j �M������R�M ��������0u�E��M�l�����Mڅ�t�U��0�Eԃ��EԹ   k��D܉E���E��M�6����MQ�UR�"���������tFj �M������Q�M �>����E��Uۃ�0|$�Eۃ�9�MԊUۈ�E�;E�s	�Mԃ��M���Uڅ�u�E܉EԋM�� �E�    �U�Rj
�E�P�M�Q��������E��E�    �UR�EP�[������ȅ�t	�UЃ��UЍE�9E�t�}� u�M�;M|�U;U�}�EЃ��E���M�Ủ�EЋM�3��������]����������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��  ���3ŉE�VP�E�d�    ������ǅ|���    h�  h��E�HQ�R�E�HQ�R������E��tQ������Q�M����������������������E�    �����P�e�������p����E������������I����O������Q�M�W����������������������E�   ������P�1�������p����E����������������ƅ���� ƅw��� �M��\���E�   ��D���Q��p��������M��;���E�������R�M������������������������E�������Q�F�������4����E��������t����UR�   k�����Q�   k� ��P��4�������ǅX���    ���X�������X������������D  ��X����7  ��X�����D�����L�����L����� ��L�����L���X�  ��L������v�$��v�U�R��p���������E������������E��M�F����u=�EP�MQ�C������Ѕ�t&�M�������M������� ;�tj �M��{����Q��X���uH�M��������w;�MQ�UR�����������u�M�g������M������;�t
j �M��(�����x���R�M������������������������E�������Q������s����E���x����<����������d����M�n����UR�EP�Z������ȅ�tv��l���R�M����������������������E���|�������|���������R�������������t)�M����������������;�uǅ8���   �
ǅ8���    ��8�����_����E�   ��|�����t��|������l����`�����_�����t������T���R�M�������������������������E�	������Q������տ����T����E���T���������T�����tƅ�����E������������E��M�������  �EP�MQ��������Ѕ�t�t  ������P��p����<����������������� ����E�
��|�������|����� ����y�����vej ������P��p���������������������������E�   ��|�������|���������������0�M�������;�uǅ$���   �
ǅ$���    ��$�����g����E�
   ��|�����t��|����������������E�   ��|�����t��|�����������������g�����t?�M����������R��p���� ���������������P�M��N��������������!  ��,���Q��p���誼���������������������E���|�������|����������&�����vej �����Q��p����b����������������������E�   ��|�������|���������蟿���0�M������;�uǅ(���   �
ǅ(���    ��(�����f����E�   ��|�����t��|�����������E�   ��|�����t��|������,����|�����f�����tF�M莾��������P��p���莻��������������Q�M�������������7���ƅw�����   ������R��p��������������������������uǅ0���   �
ǅ0���    ��0�����U����������������U�����t�f��H���R��p�������������������������uǅ<���   �
ǅ<���    ��<�����W�����H����v�����W�����tƅw�����  ǅ`���    ��p����E�����H�����d���R��p��������E���d���������u	ƅo��� ���p����V�����o�����o�����n�����n�����t��d����н�����|e��M������EP�MQ��������Ѕ�t?�M�Y�����P�MQ�v�������h�����h���
s��h�������P�M�覽����L  j j�M������E�ǅx���    ��M�w����MQ�UR�c�����������   �M�������Q�UR���������h�����h���
sV��h�������Q�M��#�����x���R�M�蒼��� ��t'��x���Q�M��{�����,�����,������,�����K��x���R�M��R���� ��t�M�C�������n���;�t�"�j j�M�������x�������x���������x��� u�.��x���Q�M���������~��x�������x����ƅ������d���������P�������������   ��x��� ��   ��P������u
�   �   ��x�������x���t��P����2��x���P�M��j����;�u(��x��� u(��P����2��x���P�M��B����;�}	ƅ�����%�   �� ��P������~��P�������P����A�����������t �E��M��J����E���d����;�����  �E��M��*�����p����ҽ����l����MQ�UR�*�����������   ��l�������   �M��������l���;���   �MQ�M����P��������Ѕ�t\��`���;�H���}N�M�J�����Q�UR�g�������h�����h���
s'��h�������Q�M�藺����`�������`���눋�`���;�H���}ƅ�����M��#�����u	ƅ�����+���`�������`�����`���;�H���}j0�M��3������E���d���������   ��X���u�vƅm��� ��M������EP�MQ��������Ѕ�t)�M�`�����PjH��4����o����ȅ�t	ƅm���븋�X�����D����� u��m�����uƅ������������������  �M��:�������  �����������E���<���P�M������������������������E�������R����������E���<����������M������`���P�M��K����������������������E���|����� ��|���������P�����輿�����<����ȅ�t@�UR�EP�������ȅ�t)�M�#���������������;�uǅ@���   �
ǅ@���    ��@�����e����E�   ��|����� t��|���ߍ�`����������e�����t������H���P�M��m����������������������E�������R������t�����V����E���H���������V�����tƅ�����E������蓵����������tj �M��������w�����tj-jj �M������E�P�M�������|�����@��|����E��M��M����E������M��>����E�M�d�    Y^�M�3��������]� ��sEi�kGo3t  �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��E�    ����P�M�����E����E��E��]� ����������������U��j�h�d�    PQ��@���3ŉE�SVWP�E�d�    �e��M��E�P�M�;����}���,�   ���M�����E��M��A    �U��B    �E��@    �M��A    �E�    �U���,Rj �E��HQ�¶�����E��U��E��B�M�Qj �M��������M�����j j �����|��E�������E������U��B(��t�M��Q(�U��	�E��H)�M��U��E��P�M��y |	�U��z|
�E��@    �M��Q.R�E��H*Q�U��B+P�M��� Q�M�������U��B/P�M��Q,R�E��H-Q�U���$R�M������E��t,jhȦ�M��� Q�,�����jhȦ�U���$R�������M�d�    Y_^[�M�3��|�����]� �������������������������������������������������������������������������������������������������������������������������U����M��E�P�M������P�E��H�P��]� �����������������������U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��j�h�d�    PQ��SVW���3�P�E�d�    �e��M�E��@    �M��A    �U��B    �E�    �EPj �M�������M�����E�M�U�Q��M������j j �;����x~��E�������E������M�d�    Y_^[��]� ���������������������������������������������U��j�h�d�    P�����3�P�E�d�    �M�E�P�M������E��M��M��E�    �U�R�M��讲���E������M�������M�d�    Y��]� �����������������������������U��j�h�d�    P��   ���3�P�E�d�    j j ��������   ������#Uu�   �} um�@����E�j'hа�E�Pj�õ�����E��E�    �}� tj �MQ�M������E���E�    �U�U��E������P��,���P�E�P�M�)���� �P�����P�MQ������P�M����j j �ӫ�����   ������#Uu�   �} um�����E�j(hа�E�Pj�������E��E�   �}� tj �MQ�M������E���E�    �U�U��E������T��x���P�E�P�M�u���� �T��_���P�MQ�˾����P�M�S���j j �q������   ������#Uu�   �} um������E�j)hа�E�Pj�[������E��E�   �}� tj �MQ�M��H����E���E�    �U܉U��E������X��Ĭ��P�E�P�M������ �X�諬��P�MQ�F�����P�M蟻��j j �"������   ������#Uu�   �} um�$����E�j*hа�E�Pj觳�����E��E�   �}� tj �MQ�M��e����E���E�    �UԉU��E������\�����P�E�P�M����� �\������P�MQ������P�M����j j ��������   ������#Uu�   �} uo�p����E�j+hа�E�PjX�������E��E�   �}� tj j �MQ�M��5����E���E�    �ỦU��E������`��Z���P�E�P�M�W���� �`��A���P�MQ�>�����P�M�5���j j �������   ������#Uu�   �} uo�����E�j,hа�E�PjX�=������E��E�   �}� tj j �MQ�M������E���E�    �UĉU��E������d�褪��P�E�P�M衹��� �d�苪��P�MQ�k�����P�M����j j �6������   ������#Uu�   �} us�����E�j-hа�E�PjD臱�����E��E�   �}� tj �MQ�M��-����E���E�    �U���|����E������h�����P��|���P�M����� �h��ѩ��P�MQ�!�����P�M�Ÿ��j j ��������   ������#Uu�   �} uy�J�����x���j.hа��x���Pj�ǰ�����E��E�   �}� tj �MQ�M��Z����E���E�    �U���t����E������l��-���P��t���P�M�'���� �l�����P�MQ�������P�M�����M�d�    Y��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��E��H(��u,�}w&�}w �}wkU�E��kU(��x��E���E�Ȧ�M��M�j�U�Rj�EP芪������]� �������������������������U��j�hPd�    P�����3�P�E�d�    �E�   �} u	�E�    ��EP�M蝵���E��M��M��E� �M������E������M�����E�M�d�    Y��]������������������������������������U��j�h�d�    P���3�P�E�d�    �E�    ��E ���E �M躙���M蕬���}  v�M�$������R�M��������_����E�M��U�P�E������M�/����E�M�d�    Y��]�����������������������������������������U��j�hId�    P��  ���3ŉE�P�E�d�    ��X����E�    h  h��EP�,������M��tK������R�M�,����������������������E�������Q���������8����E� �������Ә���I��t���R�M������������������|����E���|���Q辻������8����E� ��t���舘���U�R��8����]����E���8������������������ }������؉����������������������@����M$袭��;�@���w(�E@P�M$荭����@���+ȃ�Qj �M$�������   �M��t��������   �M��`���� ����   ��8���������/����M��<�����0����M$�$���+�@�����(�����0������tx��0������~k��0����;�(���sZ��0������(���+�(�����/���Qj��(���R�M$�����   �� ��0������~��0�������0����z����M������E��M ��tH��`���R��8����ͯ��� ������M�Q��8���詞����x�����x���R�M������M��U����L��H���P��8����B�����������H���R��8�������������������P�M��������H��������M�������E��M������t2��d���Q��8����^���������������R�M�������d���輧��ƅ?��� ǅD���    ǅ4���    ���4�������4�����4����  ��4����������$�����$����� ��$�����$���X��   ��$��������$����M������D�����D����   �M������D�����D����   ��@��� vǅ���   �
ǅ���    �M$�ɪ��;�@���w�M$蹪����@���+ȃ�������
ǅ���    �M$蔪�����������D�����D������D�������D�����4���tƅ?���������M���������������������� |1	������ v&�M����;�D���v�M����+�D���������
ǅ���    �������D����M����%�  ����������@tO�����   u��?�����u8��D���R�EP�MQ�UR������P许������P�M�UǅD���    ǅ4���    ���4�������4�����4����  ��4���������� ����� ����� �� ����� ���X��  �� �������$����M�����P�����P�M������������������������E����̉�@���������R�b�����8����EP�MQ������R��������������������P�M�U�E������莲���5  �M�膨������   j��$���P�M������������������������E����̉�0���������R�������L����EP�MQ������R���������������������P�M�U�E���$���������  ��@��� ��   �M$����P�����P�M$�i����������������������E����̉�P���������R�2�����p����EP�MQ������R�`�������������������P�M�U�E�������^����  �M$�V���;�@����	  �E@Pj �M���������������J�����8���������Qj �M��������������#����M$�������@���+�R�E@P�MQ�UR��|���P��������P�M�U�M$�Ʀ��P������P�M$�L����������������������E�	���̉�d���������R������<����EP�MQ��l���R�C�������������������P�M�U�E��������A����y  �M$�9���+�@���P������P�M$�����������������������E�
���̉�\���������R������D����EP�MQ��t���R谽������������������P�M�U�E�������讯����8����x�����Pj �M�W������5�����������@���Q��@���R������P������Q�M$�����������������������E�������膢���������������������E����̉�T���������R������4����EP�MQ������R�Լ������������������P�M�U�E��������Ү���E��������î���mj�EP�MQ�UR������P躳������P�M�U�����   u8��D���P�MQ�UR�EP������Q耳������@�U�EǅD���    ������M��L�������   �M��;�����Pj�� ���Q������R�M������������������� ����E��� ����p����������������������E����̉�l���������R�]�����h����EP�MQ������R苻������������������P�M�U�E��� ���艭���E��������z���j j �M�ʡ����D���P�MQ�UR�EP�MQ�e������E��M��d����E��M��X����E� �M��L����E������M$�=����E�M�d�    Y�M�3�������]�< ��g������.� �I Òn������0� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E���E�M� ����} v�MQ�M�b�����������ӋU�E��M�J�E]����������������������������U��Q�M��E��HQ�0������U��BP�!������M��QR�������E��HQ��������]��������������������������U��Q�M��E��HQ�Ч�����U��BP��������M��QR貧������]�������������������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M���]� ���U����M�j_hP��EP�MQ觩����j`hP��UR�EP萩�����M���Q�UR�EP�MQ�UR��������E��}� }	�E�������}� u	�E�    ��E�   �E��E�E��]� �����������������������������������U����M��E�    �E��HQ�M������U����U��E��]� ���������������U��Q�M��E��@��]����������������U��Q�M��E��@��]����������������U��Q�M��E��@��]����������������U����M��E�    �EP�M跞���M����M��E��]� ������������������U��j�h�d�    P��D���3ŉE�P�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M������E�    �EP�MQ�e������Ѕ�t�E$����U$�
�M��:�����u�E$����U$�
�P�M��)����E��E�    �E�Pj �M�Q�U�R�)������]��E�;E�t�}� t�M$����E$���M(�E���U�E��M�J�E������M��ז���E�M�d�    Y�M�3�膧����]�$ �����������������������������������������������������������������������������������U��j�h�d�    P��<���3ŉE�VP�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M��u����E�    �M������E��EP�MQ�������Ѕ�t�E$����U$�
�}� u�E$����U$�
�   �E�    �E�P�M(�W���j �M��U������-u)�UĉU��E�P�M(�;����   k�
�L��Uă��U��	�Eă��EċM�;M�s#�U�R�M������0�E�P�M(������L5���̋U�E��M�J�E������M��*����E�M�d�    Y^�M�3��إ����]�$ �����������������������������������������������������������������������������������������������������U��j�h8d�    P��p���3�P�E�d�    �M��E�P�M������E܋M܉M��E�    �U�R�������E��E������M�谂���E�    �E(�E�M��A�M�}�8�K  �U������$�$��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�辰����P�M�U�  �E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�������@�U�E��  h(��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�������P�M�U�  �E�P�M�Qjcj �UR�EP�M�Q�v������U �M ��U ���ukM�d��l  �U$�J�Q  �E�P�M$��Qjj�UR�EP�M�Q�*������U �M ��  hD��U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��I����P�M�U��  �E�P�M$��Qjj �UR�EP�M�Q�������U �M ��  �U�R�E$��Pjj �MQ�UR�E�P�������M �U ��~  �E�P�M$��Qhn  j�UR�EP�M�Q�T������U �M ��I  �U�R�E�Pjj�MQ�UR�E�P�%������M �U ��E ���u�U���E$�P�  �M�Q�U$��Rj;j �EP�MQ�U�R��������M �U ���  hT��E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M���}����@�U�E�  hX�j �MQ�UR踎�����E�}� }�E ����U �
�kE��M$A�U$�B�Q  hh��E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��{}����@�U�E�  h|��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��>}����P�M�U��  �E�P�M$Qj;j �UR�EP�M�Q�������U �M ��  h���U$R�E P�MQ�UR�EP�MQ�UR�E�P�M���|����P�M�U�k  �E�P�M$��Qj5j �UR�EP�M�Q�D������U �M ��9  �U�R�E$��Pjj �MQ�UR�E�P�������M �U ��  �E�P�M$��Qj5j �UR�EP�M�Q��������U �M ���   h���U$R�E P�MQ�UR�EP�MQ�UR�E�P�M���{����P�M�U�   �E�P�M�Qjcj �UR�EP�M�Q�t������U �M ��U ���u �}�E}�M��d�M���U�U��E$�M��H�B�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��o�����P�M�U��E ����U �
�EP�MQ譤�����Ѕ�t�E ����U �
�E�M��U�P�E�M�d�    Y��]�( �I ��̟A�����+�סǢ�3�p�ԣ�����]���	�F������C�Τ 	
	 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hhd�    P��D���3�P�E�d�    �M�h  h���EP�MQ�UR�EP�O�����h  h���M$Q��������U�R�M�U����E��E��E��E�    �M�Q�ל�����E��E������M��z���M��Q����E�}� u�E�   �UR�EP�f������ȅ�t�  �M������Rj�M���������u?�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��}�����P�M�U�E�   �   �}�u>�E�P�M$��Qjj�UR�EP�M�Q�������U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P�л�����M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��������@�U�E�MQ�UR�q���������t'�M������QjH�M�������Ѕ�t
�M�I����EP�MQ�3������Ѕ�t<j �M訒����P�M��O����E��M��:t�U��,t	�E��/u�M�����MQ�UR�����������t'�M�W�����QjH�M��i����Ѕ�t
�M踂���EP�MQ�s������Ѕ�t��   �M������Pj�M��&����ȅ�uW�}�u�U ����M ��@�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��u�����P�M�U�}�u�E�   �w�}�t�}�u>�E�P�M$��Qjj�UR�EP�M�Q�������U �M ��U$�B���M$�A�-�U�R�E$��Pjj�MQ�UR�E�P�Ź�����M �U ��EP�MQ蛗�����Ѕ�t'�M������PjH�M��$����ȅ�t
�M�s����UR�EP�]������ȅ�t<j �M�Ґ����R�M��y����E��E��:t�M��,t	�U��/u�M�����EP�MQ�
������Ѕ�t'�M聐����PjH�M�蓧���ȅ�t
�M�����UR�EP蝝�����ȅ�t�U ����M ��  �M�1�����Rj�M��C�������uM�}�t�M ����E ��3�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�蒠����P�M�U�   �}�u>�E�P�M$��Qjj�UR�EP�M�Q�0������U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P�������M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�������@�U�E�MQ�UR�^���������t�M ����E ��M�U��E�A�E�M�d�    Y��]�  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M�h}  h���EP�MQ�UR�EP������h~  h���M$Q�|������U��BPj �MQ�UR�ˁ�����E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U��j�h�d�    P�����3�P�E�d�    �M�h�   h���EP�MQ�UR�EP������h�   h���M$Q�������U�R�M�����E�E�E��E�    �M�Q藔�����E��E������M���q���U�R�E$��Pjj �MQ�UR�E�P�j������M �U ��E �8 uj �M�ċ����Q�M��k����Ѓ�:t�E ����U �
�2�E�P�M$��Qj;j �UR�M�|��P�E�P�������M �U ��E �8 uj �M�]�����Q�M������Ѓ�:t�E ����U �
�/�E�P�M$Qj;j �UR�M�{��P�E�P蟳�����M �U ��E�M��U�P�E�M�d�    Y��]�  ����������������������������������������������������������������������������������������������������������������������������U����M�hn  h���EP�MQ�UR�EP�������ho  h���M$Q茾�����U��BPj �MQ�UR��~�����E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U��j�h�d�    P�����3�P�E�d�    �M�h�  h���EP�MQ�UR�EP������h�  h���M$Q譽�����U�R�M�%����E�E�E��E�    �M�Q觑�����E��E������M���n���E�    �U�R�E�Ph�  j �MQ�UR�E�P�s������M �U ��E ���u6�}�l  |�U���l  �U���}��   ~�E ����U �
�E$�M��H�U�E��M�J�E�M�d�    Y��]�  ��������������������������������������������������������������������������������U����M��E�    �E��HQ�M諳���U����U��E��]� ���������������U��Q�M�j{hP��EP�MQ艏�����U+UR�EP�ը������]� �������������������������U��Q�M��E��H$�U�
�E��]� ���������������������U����M��E�    �E��HQ�M�����U����U��E��]� ���������������U��Q�M������]� ����������������U��Q�M��E��H �U�
�E��]� ���������������������U����M��E�    �E��HQ�M�[����U����U��E��]� ���������������U��j�h d�    P��X���3ŉE�P�E�d�    �M��E�P�M�J����E��M��M��E�    �U�R�̎�����E��E������M���k���E�P�   k���l�R�   k� ��l�Q�M������E� �E�    �M �H����Ѕ�u+j �M �Mx��� �   k�
�L�;�u�E��U����U��M ������E��E��E��	�M����M��U�;U�s%�E�P�M ��w�����R�E�P贒������
s�ʋM�+M�Q�U�R�M ��w��P�M�耖���E�   �M�袺������t�   k� �D�Pj�M�葄���   k� �D�P���̉e��U�R�-����E��E�P�MQ�UR�EP�MQ�UR�EP�M�胙���E������M��7|���E�M�d�    Y�M�3�������]� �����������������������������������������������������������������������������������������������������������������������������������U��j�hPd�    P��p���3ŉE�P�E�d�    �M��E� ���] ����Au�E��E ���] �E�    �	�E���
�E��E ������u�}��  s�E �5���] �Ѓ��E �$h�j(�M�Q�&������E��}� }�U�E��M�J�E��   �U�R�M�Z����E��E��E��E�    �M�Q�܋�����E��E������M��i��j0�M�螴���E�j �U�R�M��"���E�   j �M��t��P�E��L�Q�   k� �L�Q�M������U�R�E�P�M��H����M�Q���̉e��U�R�����E��E�P�MQ�UR�EP�MQ�UR�EP�M��C����E������M���y���E�M�d�    Y�M�3�覊����]�  �������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��P���3ŉE�P�E�d�    �M�h  h���EP虞����h	  h���MQ�M������|��U蠀��E�M��ܵ���E�    �M$��u�   ��E �D���   ��U$�T�   k��U �T��E�   ��E����E�j �M�Q�M�蝀���M��������P�UR�E�P�M��b|��P�M�Q�M������E��U��U��E��M�����P�������E��}� v	�E�   ��E�    �E��E��E� �M������M˅�t��i����UR�EP�M�Q�M��q��Pj�M��q��P�UR�������E������M���w���E�M�d�    Y�M�3�莈����]�  �����������������������������������������������������������������������������������������������������������U��Q�M��E��@��]����������������U��j�h�d�    P��\���3ŉE�VP�E�d�    �M��E�    jhhP��EP�MQ�M������M��ʳ���E�    �U+U�Ũ}� ��   �E�P�M��]����M���Q�UR�EP�M�Q�M������E��U��U��E��M��5������M��gz���V�E�P�M������E��M��M��E��M�����P�4������E̍M��/z��9E�w	�E�   ��E�    �UȈU��E��M������E� �M�������EӅ�t��6����M�Q�M�蝩���U�R�M�u���Eă��E��E������M���u���E�M�d�    Y^�M�3�舆����]� �����������������������������������������������������������������������������������������������������U��Q�M��E�P�M�脉���M�AP�M�~����E��]� ���������������������U��Q�M��E���M��B$�Ћ�]���������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P �ҋE��]�  �������������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��EP�MQ�U���M��P(�ҋ�]� ������������U��Q�M��EP�M���M��B,�ЋE��]� ���������������U����M��E�    �EP�M���M��B �ЋM����M��E��]� �������������U��Q�M��EP�M���M��B(�ЋE��]� ���������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E��H;Mr�M�}v��;Es�M��<����U��B+E;Es�M��Q+U�U�M�Nv��+E�E��E�;Es�M��M���+U�E��H+M;�w�M������U��B+E+E�E��M��QU+U�U�E��H;M�sj �U�R�M��Ck���E�;EtS�M�Q�M��2���EEP�M��#���EEP�*n�����UR�M�ٌ��EP�M������EP�Ǔ�����  �E;EwS�MQ�M��ׅ��EP�M��˅��EP��m�����U�R�M�賅��EEP�M�褅��EEP�m�����9  �E;EwS�M�Q�M��|���EEP�M��m���EEP�tm�����UR�M��R���EP�M��F���EP�Pm������   �EE;EwX�M�Q�M�����EEP�M�����EEP�m�����UR�M������MM+M�P�M������EP��l�����{�UR�M��Ƅ��EP�M�躄��EP��l�����E�P�M�袄��EEP�M�蓄��EEP�l�����M+MQ�M��u���EEP�M��f���EEP�ml�����U�R�M��m���E���]� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��} th�  h ��EP�"q�����MQ�M���[���Ѕ�t+�EP�M��C����M+�Q�U�R�EP�MQ�M��v���  �U��B;Es�M������M��Q+U;Us�E��H+M�M���+U�E��H+M;�w�M��~����U��B+E+E�E��M;Ms*�U�R�M�蹂��EEP�M�誂��EEP�j�����} w�} v~�E��HM+M�M�j �U�R�M��og������tZ�M;Ms*�U�R�M��W���EEP�M��H���EEP�Oj�����EP�MQ�M��)���EP�������U�R�M���j���E���]� �������������������������������������������������������������������������������������������������U��j�h�d�    P��   ���3�P�E�d�    �M��E�   �E,P�M �C����ȅ���   ���̉e��UR�{����EȋEȉE��E����̉e��UR�]����E��E��������EЋE�P��p���Q�M��B����E��U��U��E����̉e��E�P�����E؋M؉M��E����̉e��UR������E��E�讙�����E�E�P�M������E���p����>z����   �M Q�M,�q���P�M ����P���̉�|����UR蠎���E�E�E��E����̉e��UR肎���E��E��4������E�E�P��d���Q�M��g����E܋U܉U��E����̉e��E�P�?����E̋M̉M��E�	���̉e��UR�!����E��E��Ә�����EċE�P�M�蟫���E���d����cy���M��M��E��M�bc���E��M�Vc���E� �M �9y���E������M,�*y���E��M�d�    Y��]�0 ��������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M�j �EP�M��i����]� ���������������������U��Q�M��E��M;Hw�UR�M��[g����EP�M��U+QR�M��Ar����]� �������������������U��Q�M��E���M��B�Ћ�]���������U��j �EP�MQ�UR��}����]����������������������U���   ���3ŉE��E��\����MQ�UR�Ԉ�����E��E�����X����} t	�M�    �U�����U��}��  j��l���P�MQ�UR��\���P跆������h���Q�h��$j�M�Q�EX������h��� uQ���$j�U�R�(X�����   ǅx���   �   �� ��l���Qj�U�R��W������x���;�h���}Y�M�Qj�U�Rj�E�P�[������x�������x�����x������l���Pj�M�Q�W����j�U�Rj�E�P�W����뙋MQ�   k� �M�l���Q�U�R蘊����ٝ|����d  �}��*  j��l���P�MQ�UR��\���P�+�������`���Q�d��$j�M�Q�W������`��� uQ���$j�U�R�W�����   ǅt���   �   �� ��l���Qj�U�R�V������t���;�`���}Y�M�Qj�U�Rj�E�P�Z������t�������t�����t������l���Pj�M�Q�[V����j�U�Rj�E�P�tV����뙋MQ�UR�E�P耉����ٝ|����   k� ��l���P��|���Q脈�����0�}�u��ٝ|�����}�u��ٝ|������ٝ|�����X��� t-��|���R��g������d�����d������ �  ��d���f�
م|����M�3��yw����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�y����]����������������������U���(  ���3ŉE��E�������MQ�UR褄�������������������������} t	�M�    ����������������������  j�E�P�MQ�UR������P�{�����������������$j�M�Q蓁���������� u�����$j�U�R�t������   ǅ����   �   �� �L�Qj�U�R������������;�����}Y��0���Qj�U�Rj�E�P���������������������������D��Pj�M�Q萀����j�U�Rj�E�P�@�����뙋MQ�   k� �ML�Q�U�R������ݝ�����t  �������1  j�E�P�MQ�UR������P���������������p��$j��`���Q�k����������� u�����$j�U�R�L������   ǅ����   �   �� �L�Qj�U�R�����������;�����}b�� ���Qj��`���Rj�E�P��������������������������D��Pj��x���Q�b����j��x���Rj�E�P������됋MQ�UR�E�P�������ݝ�����   k� �D�P������Q�,������6������u�h�ݝ�����������u�x�ݝ�������ݝ���������� t-������R�s������������������� �  ������f�
݅�����M�3��/s����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�z����]����������������������U���(  ���3ŉE��E�������MQ�UR�T��������������������������} t	�M�    ����������������������  j�E�P�MQ�UR������P�+~����������������$j�M�Q�.����������� u�����$j�U�R�������   ǅ����   �   �� �L�Qj�U�R苂����������;�����}Y��0���Qj�U�Rj�E�P訂�������������������������D��Pj�M�Q�:�����j�U�Rj�E�P������뙋MQ�   k� �ML�Q�U�R�D�����ݝ�����t  �������1  j�E�P�MQ�UR������P衛�������������p��$j��`���Q������������ u�����$j�U�R�������   ǅ����   �   �� �L�Qj�U�R�c�����������;�����}b�� ���Qj��`���Rj�E�P�}��������������������������D��Pj��x���Q������j��x���Rj�E�P踁����됋MQ�UR�E�P������ݝ�����   k� �D�P������Q������6������u��ݝ�����������u���ݝ�������ݝ���������� t-������R�d������������������� �  ������f�
݅�����M�3���n����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} u�E�E�M�M��	�U����U��E��Q���������t��U����-t�M����+t	�E�+   ��E���M��U����U��E��E��MQ�UR�EP�M�Q��{�����E�U�E�;u�M�U��E�M;u�}� u$�U���+u	�}����w�E���-uC�}�   �v:�Ĕ��� "   �} t	�M�   �U���-u	�E�   ���E�����E����E���-u
3�+M�M���U�U�E��]���������������������������������������������������������������������������������������U��j �EP�MQ�UR��z����]����������������������U���$�} t	�E�     �M�M��	�U����U��E��Q�L�������t��U����-t�M����+t	�E�+   ��E���M��U����U��E��E��} |�}t�}$~�} t�M�U�3���  �   �} ~D�}u<�E����0u1�   �� �E����xt�   �� �E����Xu	�U����U��U�E����0t	�E
   �A�   �� �E����xt�   �� �E����Xu�E   �U����U���E   �E��E��	�M����M��U����0u���E�    �M��M��E�    �	�U����U��EP�M��R�Z�����P�   k� ����Q�,q�����E�}� t#�U�U�E�-���E��M��M�U�ʉM�렋E�;E�u�} t�M�U�3��   �E�+E܋M����+E�y�L�}� !�E��M�+�9M�r�U��E�+�3��u;E�t%趑��� "   �} t	�E�    �E������E�+�M���-u3�+U�U�} t�E�M���E��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�|w����]����������������������U���(�} u�E��E�M�M��	�U����U��E��Q���������t��U����-t�M����+t	�E�+   ��E���M�U����U��E�E��MQ�UR�EP�M�Q跓�����E�U�U�E�;u�M�U��E�M;u�U�U�u4�E���+u�}����w"r�}��w�M���-u\�}�   �rSw�}� vK诏��� "   �} t	�U�   �E���-u�E�    �E�   ���E������E�����E��U��2�0�M���-u3�+U�    E�U؉E���M�M؋U�U܋E؋U܋�]���������������������������������������������������������������������������������������������U��j �EP�MQ�UR�e�����]����������������������U���<V�} t	�E�     �M�M��	�U����U��E��Q��������t��U����-t�M����+t	�E�+   ��E���M�U����U��E�E��} |�}t�}$~�} t�M�U�3�3��]  �   �} ~D�}u<�E����0u1�   �� �E����xt�   �� �E����Xu	�U����U��U�E����0t	�E
   �A�   �� �E����xt�   �� �E����Xu�E   �U����U���E   �E��E��	�M����M��U����0u���E�    �E�    �M��M��E�    �E�    �E� �	�U����U��EP�M��R������P�   k� ���Q��k�����E��}� t@�U܉UԋE��E؋M�����M��E�RP�U�R�E�P�i����ȋ��E����M܉u�냋U�;U�u�} t�E�M�3�3���   �U�+U�E���+щU�y�   �}� Y�E���M�+ȋE�M̉EЋM�;M�r<w�U�;U�r2�E���M�+ȋu��E�RPVQ�]���EĉUȋU�;U�u�E�;E�t,����� "   �} t	�M�   �E������E������E�+�U���-u3�+Eܹ    M��E܉M��} t�U�E���E܋U�^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����i���E���D���   �� ��U��}� t�E�P��r�����E��E��U���]�����������������U���$�E�    �E+E�E�M+M�M��} u�D���   �� ��E��h���E���M�Q�U��E��M܃}� ui�U�;U�}�E�E���M��M�U�R�EP�MQ��L�����E�}� u(�U�;U�t �E�;E�}	�E�������E�   �M�M���U�U��E��E��M�M�Q�U�R�EP�M�Q�URh   �E�Pj �hk���� �E��}� u袉���    �E�����	�M����M��E���]���������������������������������������������������������������������������U���3�f�E�3�f�M�j�U�Rj"�BC���   k��P�@�����   k� �D���0u	�E�   �I�   k� �D���1u	�E�   �(�   k� �D���2u	�E�   ��E�    �M��M�U�U��E���]���������������������������������������������������U���l���3ŉE�VW�} t�} u3��@  �E���u�} t3ҋEf�3��!  �} u�M�Q�~�����   ���}��UЉU�E�x t�} t�Mf��Ef��   ��  �M�yt,�U�zt#hH�hpjj j^h��j�FA������u̋M�9 ��   �   �� �E�M�	��U�zv6�} t	�E�   ��E�    �E�P�MQj�URj	�E�Q���u�U�    �:���� *   ����(  �E�     �M�A�  �U��E��M����U�D
�Mσ��   ��#���   �E�M;Hs�   k� �M�U��������   �h�E�xv;�} t	�E�   ��E�    �M�Q�UR�E�HQ�URj	�E�Q���u$�U�B��u�M�    �d���� *   ����U�U�B�M�K�} t	�E�   ��E�    �E�P�MQj�URj	�E�Q���u����� *   �����   _^�M�3��\^����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��� �E+E���E�M+M���M��E�    �} u�C?���   �� ��E��	�M�Q�U��}� ui�E�;E�}�M�M���U��U�E�P�MQ�UR��   ���E�}� u(�E�;E�t �M�;M�}	�E�������E�   �U�U���E�E��M��M��G�U�R�EP�M�Q�URh   �E�P��f�����E��}� u�d����    �E�����	�M����M��E���]�����������������������������������������������������������������������������U��Q��E���E�M���M�U���U�} ~7�E��U�;�t%�M��E�;�}	�E�������E�   �E���3���]�����������������������������U����E+E���E�M+M���M��E������E�    �} u�l=���   �� ��E��	�M�Q�U�}� u)�E�;E�w�M���Q�UR�EP��E�����M�M��   jgh�j�U�R�8�����E��}� ��   �E�P�M�Q�U�R�EPh   �M�Q�sv�����E��}� u/j j �U�R�EPh   �M�Q�Mv�����E��}� u�E�����0�E�    �	�U����U��E�;E�s�M�M�f��E��Mf�A�ك}� tj�U�R�}J�����E���]����������������������������������������������������������������������������������������������U����E�Pj�MQj���u	�E�    ��U��U�f�E���]�����������������������������U��EP�M+M��Q�URj��E]����������������U��Qf�Ef�E��M����  u�_�U�z u*�E=   }�M��A|�U��Z�E�� f�E��,j�M�Qj�URh   �E�HQ�t������uf�Uf�U�f�E���]������������������������������������������������U��Qf�Ef�E��M����  u�_�U�z u*�E=   }�M��a|�U��z�E�� f�E��,j�M�Qj�URh   �E�HQ��s������uf�Uf�U�f�E���]������������������������������������������������U����E+E�E�M+M�M��E������} u��9���   �� ��E���]���E���M�Q�U�E��M��}� u*�}� u$�U�;U�w�E�P�MQ�UR�dB�����E��E��ej�M�Qj j �U�R�EPh   �M�Qj ��q����$�E��}� t7�U��U�E�;E�)j�M�Q�U�R�EP�M�Q�URh   �E�Pj �q����$�E��]������������������������������������������������������������������U����E��M��E�    �	�U����U��E��Q�2q������t��U����-u�E�   �M����M���U����+u	�M����M��U����nt�M����N��   �E����E��M����at�E����Au�U����U��E����nt�U����Nt�M��U��E�    �d�E����E��M��M��E�   �U����(uC�M����M��U��P萄������u�M����_u�׋E����)u�U����U��E��E��} t�M�U����  �E����it�U����I�"  �M����M��U����nt�M����Nu�E����E��M����ft�E����Ft�U��E��E�    �   �M����M��U��U��E���E�M����it�E����I��   �U����U��E����nt�U����Nul�M����M��U����it�M����IuM�E����E��M����tt�E����Tu.�U����U��E����yt�U����Yu�M����M��U��U��} t�E�M���   �U����0uw�   �� �U��
��xt�   �� �U��
��XuO�M����M�U����.u	�M���M�U��P�|w������u�M���M���U����U��E���E��	�M���M�U�E���E��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���l���3ŉE�V�E�    kE	�E�}-~�E-   �   k� �E�    �   �� �U�
    �E�    ��E���E�E�   �M���0u���E�    ��E���E�E�   �M�R��������tD�E�;E�M���0�EȈT̋Mȃ��M���   k� �M����   k� �E�뙋M�1�G���   k� ��
;�u	�M���M�}� u>��U���U�E�   �E���0u!�   k� �M����   k� �E�����M���M�E�   �U�P�2�������tB�M�;M8�U���0�MȈD̋Uȃ��Uȸ   k� �U�
���   k� �M�뛋U;U�}I�E�E��M��T̃�|�E��Lˀ��U��LˋE�Eȹ   k� �E����   k� �U��	�Eȃ��Eȃ}� ~-�M��T˅�u!�   k� �U�
���   k� �M��ă}� u$�UȉU��Eȃ��Eȃ}�.s���p���M��D� �}� ��  �E�    �Eș�	   ���	   +E��E���	   ����u	�E�    ��E�   �U��U���E����E��M����M��U�;U�}J�E���	   ����u�Uă��UċE��L̋UċE����MċUk�
�M��T�MċU��뜋E���et�U���E��   �M�M��U���U�E���+t�U���-t	�E�+   ��M��U��E���E�M��M��E�    �E�    ��U���U�E�   �E�Q��}������t�}� ��}kU�
�E��T
ЉU����E���-u�M��ىM��   k� �M�U��   k� �E��}� u�M��M�}� u�E�    �} t�}� t�U�U���E�E��M�U���E�^�M�3���N����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���d���3ŉE�V�E�    kE�E�}#~�E#   �   k� �E�    �   �� �U�
    �E�    ��E���E�E�   �M���0u���E�    ��E���E�E�   j�M�R�   k� ��P�Q�S�����E��}� tL�U�;U �E�-P��MԊ�h��T؋Eԃ��E���   k� �E����   k� �U��{����E�0�B���   k� � �;�u	�U���U�}� u>��E���E�E�   �M���0u!�   k� �U�
���   k� �M�����U���U�E�   j�E�Q�   k� P�P��R�����E��}� tH�M�;M>�U���P��EԊ�h��L؋Uԃ��UԸ   k� �U�
���   k� �M�뀋U;U�}I�E�E��M��T؃�|�E��L׀��U��L׋E�EԹ   k� �E����   k� �U��	�Eԃ��Eԃ}� ~-�M��Tׅ�u!�   k� �U�
���   k� �M��ă}� u$�UԉU��Eԃ��Eԃ}�$s��Ik���M��D� �   k� �M����   k� �E��}� ��  �E�    �Eԙ�   ���   +E��E���   ����u	�E�    ��E�   �U��U���E����E��M����M��U�;U�}L�E���   ����u�UЃ��UЋE��L؋UЋE����MЋU�����M��T�MЋU��뚋E���pt�U���P��   �M�M��U���U�E���+t�U���-t	�E�+   ��M��U��E���E�M��M��E�    �E�    ��U���U�E�   �E�Q�9x������t�}� ��}kU�
�E��T
ЉU����E˃�-u�M��ىMĺ   k� �M�Uĸ   k� �E��}� u�M��M�}� u�E�    �} t�}� t�U�U���E�E��M�U���E�^�M�3��:I����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�E��   �� �U��
%�  =�  u?�   �� �U��
��u�   k� �E����u	�E�   ��E�   f�E��]�[�   �� �E�������u�   k� �M����t/�   �� �M����  u	�E�������E�����f�E���3���]������������������������������������������������������������U��   k� E]�����������������U��   �� E]�����������������U���(V�E�E�   �� �U��
%�  ��f�E��M����   uB�   �� �E����u�   k� �M����u	�E�   ��E�   f�E��i  �'�E���u�M�Q��g����f�E��U���~3��@  �} ~T�E���   +�;MD�   �� �E���� �  t�����]��	���]��U�E���   ��  ��  �E���;E}<�   �� �U��
%����M�M����   �� �M�f�����  �  �   �� �E���� �  f�M�   �� �E�����ɀ   �   �� �E�f��M��U�D
��E�}�|�} |0�   �� �U�f�E�f�
�   k� 3��M�f�3��  �  f�Uf�U�3�f�E��M����h�U��t	�E�   ��E�    �   k� �U��
E�f�E��   �� �   k� �U�u�f�f��   �� 3��M�f��U���f�U��E���f�E��M�����   �U��t	�E�   ��E�    �   k� �U��
�M��   +ы���E�f�E��   k� �U��
�M����   �� �U��
�M��   +����º   k� �U�f�
�   �� �M�f�f�M�f��   �� �M�f��   �� �E��M��и   �� �M�f��U�� �  �E�= �  un�   k� �E����tZ�   k� �M�f�f��f�U�   k� �U�f�E�f�
�M����  u$�   �� �E�f�f���   �� �E�f��.�   �� �U��
�M�;�u�   k� �M����u3�����^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���<V�E�]܃} u�  �E�P�M�Q�Q����f�E��U�����   �E���t �   k� UR�T����f�E��E����   k� �E�E��u�M���t6�UR�1�����0�� �  �   k� MQ�1������� �  ;�u�4j��/�����   k� �U���
�}~�   �� �M�����  �U�����  �E�   �E�    �E�;E��  �M��U���]��E�   �E�P�M�Q�	P����f�E��U���~
�|  �r  �E���u-�M��U�E���E���;E}�M��U���\��G  �=  �E��M�+��EԋU���9U���   �E��������D��   �E��E�M���M�U�;U}�E�M����������D{�ًU��9U�}�E���E���M�;Mu	�U���U��	�E���E�M�;M�}�U�E�M�u�D�����ڋU��E�E�����]�~  �M�;M�#�E��������D{�U��U��E����E��S  �M��U���E�]ЋE��M�E����E���������Dzf�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E��M����������Dz��  �U��E���]�MQ�U�R�)N�����E�+E��M�;���   �U�E�+E�+�R�MQ�n.�����U�R�EP�-O�����M��U���e�]̋E��M�E����E���������DzM�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E����E�u	�E�   �$�M��U�D���]܍E�P�M�Q�FM�����U��U��   �E���;Eu
�   �   �M��U���]�E��M��R�E�P�M����j�M��U��P�_-�����M�Q�U��E��Q�N�����E�U��E�$��]�M��M��E��������D{�E�]���U��E���]��E��]܍M�Q�U�R�L�����E����E��D����E^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}3�U��E����������D{�M��UQ���$�EP�MQ�����뼋E��]�������������������������U����} u���b  �]  �}t2�   k� �U�
��������D{�   �� �M���������Dz�   k� �M��  �  �}t�   ��E���������Dz,�   k� �   �� �M��U��]��E���   ��   �   k� �   �� �E��M��]��   ��E��]��   k��E���������D{�M�Q�I*�����E��U�����M�f��   k� �E�M�$�   �� �E�������Dz�E��E��]��E��'�%�   k� �   �� �M��E��E��]��E��]��������������������������������������������������������������������������������������������������������U����} u�  �   k� MQ�rL����f�E��U���|<�E���u�   k� �E�����M���u�   k� �M����.  �U�U��E�M���U�E�M���U�   k� �U�
�]��EP�MQ�U�R�P��������$�EP�M�Q�s�����}~�   �� �E��E��]��E������]��E�Q�$�MQ�UR�������E�   ��E����E�M�;M}~�UR�EP�M�Q�������U�R�EP�M�Q�UR�E�P�l�������$�MQ�U�R�3�����E�P�MQ�UR�EP�M�Q�;�����UR�E�P�MQ�UR�O�����r����E��]���������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}<�UR�E��M�����$�������U��E���M��U����������Dz�볋E��]��������������������������������U��E��P�MQ�UR�u!�����E]������������������U���0���3ŉE��} ��   �   k� �U�
�M�   k� �\�   k� �L�Q�I����f�E��U���|S�E���u
j�6%�����   k� �   k� �E�D���M���~�}~�   �� �E����E�  �   k� �E����E�   �E�    ��M���M�U���U�E�;E�L  �	�M���M�}�}\�U�U�;U}=�E�E�M����������D{&�U�U�E���M�M��\��U�U�E������M����\���E�   �땺   k� �D���������Dz
��   �   �E�    �   k� �D��]؍E�P�M�Q�D����j�U�R��$�����E�P�M�Q�E�����E��$�UR�EP������   k� �D��e��]��E�Q�$�EP�MQ�������U܃��U܋E�;E�}$�M܋U��D���\��E��D����������Dz��������E�M�3��4����]�����������������������������������������������������������������������������������������������������������������������������������������������������������U����} t�} u�  �   k� �U�
��������D{�   �� �M���������Dz'�   k� �MQ��$�UR�EP�1������   �M�M�U�E���M��UR�EP�M�Q�������   k� �MQ��$�UR�EP�������E�   �	�M����M��U�;U}_�E��M����������D{K�U�R�EP�M�Q�f�����U��EQ���$�MQ�U�R������EP�M�Q�UR�EP�����됋E��]�����������������������������������������������������������������������������������������U����E��'  ���E��E��]��E�Q�$�UR�EP���������$�MQ�UR�������E��'  ���U��E��]��E�Q�$�UR�EP�������E��]�������������������������������������U����E�]�} �m  �}t�E�P�M�Q��@����f�E��U���u�   k� �U�E��
�5  �E���~&�   k� �E�E���   �� �U���
�  j�E�P�!�����M�Q�U�R��A�����   k� �U�E��
�E�e��   �� �M�3���   �   �� �M��]�   �� UR�E�P�.@����j�   �� MQ� �����U�R�   �� EP�?A�����   �� �E�U�$
�   ���M��}~(�   ��E���������D{�   k��E�����}~�   ��U���
�E��]������������������������������������������������������������������������������������������������������U����} u��  �   k� MQ�B�����Ѕ�}�   k� �U�
��s����z>�   k� �U�
��s����zj�5�����   k� �U���
�P  �E�E��M�U���E��M�U����E��   k� �E��]��}~�   �� �E��U�
�]��E����$�X	 �������]��E�Q�$�EP�M�Q�#�����E�   ��U���U�E�;E��   �M�Q�UR�E�P���������$�MQ�U�R�5�����E�P�MQ�UR�EP�M�Q������U�R�EP�M�Q�UR�E�P�z��������$�MQ�U�R�=�����E�P�MQ�U�R�EP�M�Q�E�����M����U�R�EP�M�Q�UR�EP�$�����E��]�������������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}5�U��E����������D{!�M��U����Q�$�EP�MQ�$����뺋E��]�����������������������U���8���3ŉE��} t�   k� �U�
��������Dzj�EP�	������   �} ~Q����$j�M�Q��
������U�ډUh��j�E�P�������M��t�U�Rj�E�Pj�MQ������U���Uu�,�E�Pj�M�Q������U�Rj�E�Pj�M�Q�V�����j�UR�c
�����]��E���������D{&�E���������D{�����E�������Dz�S��� "   �} t�E����U�
�EȋM�3���+����]����������������������������������������������������������������������������������������U����E�E��   k��E�����  ���  ug�   k��M����uA�   ���M����u/�   �� �M����u�   k� �U��
��u	�E�   ��E�   f�E��   ��   k��E�������u8�   ��E����u&�   �� �E����u�   k� �M����t.�   k��U��
%�  u	�E�������E�����f�E���3���]������������������������������������������������������������������������������U��   k� E]�����������������U��   k�E]�����������������U���0V�E�E�   k��E�����  ��f�M��U����  ug�   k��U��
��uA�   ��U��
��u/�   �� �U��
��u�   k� �E����u	�E�   ��E�   f�E���  �'�U���u�E�P�,����f�E��M���~3���  �} ~T�U���  +�;ED�   k��E���� �  t�h����]��	�h��]ЋU�E���   �m  �h  �E���;E}=�   k��E��������U�U��ʸ   k��E�f�����%  �   �   k��E���� �  f�M�   k��M�������   k��E�f��M��U�D
��E�}�|�} |Q�   k��E�f�M�f��   ��3��M�f��   �� 3��M�f��   k� 3ɋU�f�3��}  �x  f�Ef�E�3�f�M���U���f�U��E������   �M��t	�E�   ��E�    �   k� �M��U�f�U��   �� �   k� �M�u�f�f��   ��   �� �E�u�f�f��   k��   ��U�u�f�f�
�   k�3��M�f��L����U���f�U��E����)  �M��t	�E�   ��E�    �   k� �M���E��   +���U�f�U��   k� �E���M����   �� �M���M��   +����и   k� �E�f��   �� �U��
�M����   ��U��
�M��   +����º   �� �M�f��   ��E���M����   k��E���M��   +����и   ���M�f��   k��M�f�f�M�f��   k��E�f��   k��E��M��и   k��E�f��M�� �  (�U�� �  ��   �   k� �U��
����   �   k� �E�f�f��f�M�   k� �M�f�U�f��E�%��  ��   �   �� �U�f�
f��f�E�   �� �U�f�E�f�
�M����  uX�   ��E�f�f��f�M�   ��E�f�M�f��U����  u$�   k��U�f�
f���   k��M�f��S�   k��M���E�;�u<�   ��U��
��u*�   �� �U��
��u�   k� �E����u3�����^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���PV�E�]Ѓ} u�  �E�P�M�Q�%=����f�E��U�����   �E���t �   k� UR��/����f�E��E����   k� �E�E��u�M���t6�UR�"�����0�� �  �   k� MQ��!������� �  ;�u�4j�������   k� �U�x��
�}~�   �� �M�����  �U�����  �E�   �E�    �E�;E��  �M��U���]��E�   �E�P�M�Q�<����f�E��U���~
�|  �r  �E���u-�M��U�E�ʋE���;E}�M��U���\��G  �=  �E��M�+��E؋U���9U���   �E��������D��   �E��E�M���M�U�;U}�E�M����������D{�ًU��9U�}�E���E���M�;Mu	�U���U��	�E���E�M�;M�}�U�E�M�u�D�����ڋU��E�E�����]�~  �M�;M�#�E��������D{�U��U��E����E��S  �M��U���E�]ȋE��M�E����E���������Dzf�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E��M����������Dz��  �U��E���]�MQ�U�R�6:�����E�+E��M�;���   �U�E�+E�+�R�MQ������U�R�EP�	I�����M��U���e�]��E��M�E����E���������DzM�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E����E�u	�E�   �$�M��U�D���]ЍE�P�M�Q�S9�����U��U��   �E���;Eu
�   �   �M��U���]�E��M��R�E�P�9����j�M��U��P������M�Q�U��E��Q��G�����U��E�E�$��]�M��M��E��������D{�E�]���U��E���]��E��]ЍM�Q�U�R�8�����E����E��D����E^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}5�U��E����������D{!�M��U�����$�EP�MQ�%E����뺋E��]�����������������������U���V�} u���P  �K  �}t2�   k� �U�
��������D{�   �� �M���������Dz�   k� �M��   ��   �}t�   ��E���������Dz&�   k� �   �� �M�u���   �   �   k� �   �� �U�u���]�   ���M��]��   k��M���������D{�U�R������E��E�����U�f�
�   k� �U�E��$
�   �� �M�������Dz
�E��E��!��   k� �   �� �U�
�E�M�^��]��������������������������������������������������������������������������������������������������������U����} u�  �   k� MQ��'����f�E��U���|<�E���u�   k� �E�����M���u�   k� �M�h���(  �U�U��E�M���U�E�M���U�   k� �U�
�]�EP�MQ�U�R�!C�����з�$�EP�M�Q�$�����}~�   �� �E�E���]����u���$�MQ�UR�n%�����E�   ��E����E��M�;M}~�UR�EP�M�Q�B�����U�R�EP�M�Q�UR�E�P��$�������$�MQ�U�R��A�����E�P�MQ�UR�EP�M�Q�$�����UR�E�P�MQ�UR�7B�����r����E��]���������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}<�UR�E��M�����$��������U��E�ЋM��U����������Dz�볋E��]��������������������������������U��E��P�MQ�UR�u�����E]������������������U���@���3ŉE��} ��   �   k� �U�
�M�   k� �\ܺ   k� �L�Q��$����f�E��UЅ�|S�EЃ�u
j�6�����   k� �   k� �E�D���MЅ�~�}~�   �� �E����E�  �   k� �E����E�   �E�    ��Mԃ��MԋU؃��U؋E�;E�E  �	�M؃��M؃}�}\�U�U�;U}=�E�E؋M����������D{&�U�U؋E���M�M��\�܋U�U؋E������M����\���E�   �땺   k� �D���������Dz
�   �   �E�    �   k� �D��]��E�P�M�Q�0����j�U�R������E�P�M�Q�?���E��$�UR�EP�>�����   k� �D��e����$�EP�MQ�>�����Ũ��ŰE�;E�}$�M̋U��D���\�ԋE��D����������Dz��������E�M�3������]��������������������������������������������������������������������������������������������������������������������������������������������������U����} t�} u�   �   k� �U�
��������D{�   �� �M���������Dz)�   k� �M����$�UR�EP�������   �M�M�U�E�ЉM��UR�EP�M�Q�=�����   k� �M����$�UR�EP�0�����E�   �	�M����M��U�;U}a�E��M����������D{M�U�R�EP�M�Q�C=�����U��E�����$�MQ�U�R�������EP�M�Q�UR�EP�=����뎋E��]�����������������������������������������������������������������������������������U����E�]��E����$�EP�MQ�'�����E��]���������������������U����E�]��} �  �}t�E�P�M�Q�-����f�E��U���u�   k� �U�E��
�a  �E���~&�   k� �E�E���   �� �U���
�3  j�E�P�.�����M�Q�U�R� <�����   k� �U�E��
�E�e�   �� �M��   ����   �}��   �   �� �M���������D��   �   �� �E��]�   �� MQ�U�R�,����j�   �� EP������M�Q�   �� UR�o;�����   �� �M�E�$�   ��E��}~(�   ��U�
��������D{�   k��U���
��}~�   ���M����E��]��������������������������������������������������������������������������������������������������������������������������U����} u�  �   k� MQ�B�����Ѕ�}�   k� �U���
����Au:�   k� �U���
����Auj�m������   k� �U�x��
�L  �E�E��M�U�ʉE��M�U��ʉE��   k� �E��]�}~�   �� �U�E��
�]���E��$��  ��������$�EP�M�Q�������E�   ��U���U��E�;E��   �M�Q�UR�E�P�9��������$�MQ�U�R������E�P�MQ�UR�EP�M�Q�N�����U�R�EP�M�Q�UR�E�P�2��������$�MQ�U�R�8�����E�P�MQ�U�R�EP�M�Q�������M����U�R�EP�M�Q�UR�EP�������E��]���������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}7�U��E����������D{#�M��U�������$�EP�MQ�7����븋E��]�������������������������������������U���l���3ŉE��} t�   k� �U�
��������Dzj�EP�f
������   �} ~��� ��$j�M�Q�������U�ډUh�j�E�P��6�����M��t�U�Rj�E�Pj�MQ�6�����U���Uu�,�E�Pj�M�Q�6�����U�Rj�E�Pj�M�Q� �����j�UR�	�����]��E���������D{&�E��h�������D{�h����E�������Dz�4��� "   �} t�E����U�
�E��M�3�������]��������������������������������������������������������������������������������������U��EP������]����������������U��   k� E]�����������������U��   k�E]�����������������U��EP�MQ�5����]������������U���PV�E�]Ѓ} u�  �E�P�M�Q�=����f�E��U�����   �E���t �   k� UR�����f�E��E����   k� �E�E��u�M���t6�UR������0�� �  �   k� MQ�� ������� �  ;�u�4j�"������   k� �U����
�}~�   �� �M�����  �U�����  �E�   �E�    �E�;E��  �M��U���]��E�   �E�P�M�Q�<����f�E��U���~
�|  �r  �E���u-�M��U�E�ʋE���;E}�M��U���\��G  �=  �E��M�+��E؋U���9U���   �E��������D��   �E��E�M���M�U�;U}�E�M����������D{�ًU��9U�}�E���E���M�;Mu	�U���U��	�E���E�M�;M�}�U�E�M�u�D�����ڋU��E�E�����]�~  �M�;M�#�E��������D{�U��U��E����E��S  �M��U���E�]ȋE��M�E����E���������Dzf�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E��M����������Dz��  �U��E���]�MQ�U�R�(:�����E�+E��M�;���   �U�E�+E�+�R�MQ��������U�R�EP�&�����M��U���e�]��E��M�E����E���������DzM�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E����E�u	�E�   �$�M��U�D���]ЍE�P�M�Q�E9�����U��U��   �E���;Eu
�   �   �M��U���]�E��M��R�E�P�9����j�M��U��P�������M�Q�U��E��Q������U��E�E�$��]�M��M��E��������D{�E�]���U��E���]��E��]ЍM�Q�U�R�8�����E����E��D����E^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}5�U��E����������D{!�M��U�����$�EP�MQ�'����뺋E��]�����������������������U���V�} u���P  �K  �}t2�   k� �U�
��������D{�   �� �M���������Dz�   k� �M��   ��   �}t�   ��E���������Dz&�   k� �   �� �M�u���   �   �   k� �   �� �U�u���]�   ���M��]��   k��M���������D{�U�R�7������E��E�����U�f�
�   k� �U�E��$
�   �� �M�������Dz
�E��E��!��   k� �   �� �U�
�E�M�^��]��������������������������������������������������������������������������������������������������������U����} u�  �   k� MQ�����f�E��U���|<�E���u�   k� �E�����M���u�   k� �M����(  �U�U��E�M���U�E�M���U�   k� �U�
�]�EP�MQ�U�R������з�$�EP�M�Q�������}~�   �� �E�E���]����u���$�MQ�UR������E�   ��E����E��M�;M}~�UR�EP�M�Q������U�R�EP�M�Q�UR�E�P�<�������$�MQ�U�R�������E�P�MQ�UR�EP�M�Q������UR�E�P�MQ�UR�p�����r����E��]���������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}<�UR�E��M�����$�������U��E�ЋM��U����������Dz�볋E��]��������������������������������U��E��P�MQ�UR�������E]������������������U���@���3ŉE��} ��   �   k� �U�
�M�   k� �\ܺ   k� �L�Q�����f�E��UЅ�|S�EЃ�u
j�v������   k� �   k� �E�D���MЅ�~�}~�   �� �E����E�  �   k� �E����E�   �E�    ��Mԃ��MԋU؃��U؋E�;E�E  �	�M؃��M؃}�}\�U�U�;U}=�E�E؋M����������D{&�U�U؋E���M�M��\�܋U�U؋E������M����\���E�   �땺   k� �D���������Dz
�   �   �E�    �   k� �D��]��E�P�M�Q�0����j�U�R�a������E�P�M�Q����E��$�UR�EP������   k� �D��e����$�EP�MQ������Ũ��ŰE�;E�}$�M̋U��D���\�ԋE��D����������Dz��������E�M�3��������]��������������������������������������������������������������������������������������������������������������������������������������������������U����} t�} u�   �   k� �U�
��������D{�   �� �M���������Dz)�   k� �M����$�UR�EP��������   �M�M�U�E�ЉM��UR�EP�M�Q������   k� �M����$�UR�EP�y�����E�   �	�M����M��U�;U}a�E��M����������D{M�U�R�EP�M�Q�'�����U��E�����$�MQ�U�R������EP�M�Q�UR�EP�;����뎋E��]�����������������������������������������������������������������������������������U����E�]��E����$�EP�MQ�R�����E��]���������������������U����E�]��} �  �}t�E�P�M�Q�r-����f�E��U���u�   k� �U�E��
�a  �E���~&�   k� �E�E���   �� �U���
�3  j�E�P��������M�Q�U�R�=�����   k� �U�E��
�E�e�   �� �M��   ����   �}��   �   �� �M���������D��   �   �� �E��]�   �� MQ�U�R�,����j�   �� EP�8������M�Q�   �� UR������   �� �M�E�$�   ��E��}~(�   ��U�
��������D{�   k��U���
��}~�   ���M����E��]��������������������������������������������������������������������������������������������������������������������������U����} u�  �   k� MQ�������Ѕ�}�   k� �U���
����Au:�   k� �U���
����Auj�������   k� �U����
�L  �E�E��M�U�ʉE��M�U��ʉE��   k� �E��]�}~�   �� �U�E��
�]���E��$�>�����������$�EP�M�Q������E�   ��U���U��E�;E��   �M�Q�UR�E�P���������$�MQ�U�R��	�����E�P�MQ�UR�EP�M�Q�
�����U�R�EP�M�Q�UR�E�P�
��������$�MQ�U�R�
�����E�P�MQ�U�R�EP�M�Q�K
�����M����U�R�EP�M�Q�UR�EP�*
�����E��]���������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}7�U��E����������D{#�M��U�������$�EP�MQ�	����븋E��]�������������������������������������U����E�$���  ��]�����������U���l���3ŉE��} t�   k� �U�
��������Dzj�EP�[������   �} ~��� ��$j�M�Q�������U�ډUh�j�E�P������M��t�U�Rj�E�Pj�MQ�d�����U���Uu�,�E�Pj�M�Q�x�����U�Rj�E�Pj�M�Q�.�����j�UR������]��E���������D{&�E���������D{�����E�������Dz����� "   �} t�E����U�
�E��M�3�������]��������������������������������������������������������������������������������������U���V�   �� �M��� �  f�U��   f�E��   �� �U�
���E��   �� �Uf�E�f�
�M��u�   k� �M����e  �   �� �M���u:�   k� �   �� �E�uf�f��   k� 3ɋUf��E���f�E��f�M�f��f�M��   �� �E����   }W�   �� �E���   k� �U���Ⱥ   �� �Ef��   k� �Ef�f��   k� �Uf���f�E�f��f�E��   �� �U�
=   |W�   k� �E����   �� �E���ʸ   k� �Ef��   �� �Uf�
f��   �� �Uf�
뇸   �� �M����   �� �Mf��   �� �E��M�и   �� �Mf�f�E�^��]�����������������������������������������������������������������������������������������������������������������������������������������������U��E��t���� !   ��M��t���� "   ]��������������������U����E�E��   �� �U��
%�  ��f�E��M����   uB�   �� �E����u�   k� �M����u	�E�   ��E�   f�E��Z  �1�   �� �M�������u�   k� �U��
��u3��'  �M���   +��E+�f�U��M���3��  ��   �U���|B�   �� �M���� �  �   �� �M�f��   k� 3ɋU�f�����   �   �E���f�E,�f�M�f�U�f��f�U��E���L��U��J�M�#�f�M��U���L��M��U��B3��M���L��M�f�Q�U���~*�   k� �U��
�M��f�M��   k� 3ɋU�f��E���t	�E�������E�    f�E��]��������������������������������������������������������������������������������������������������������������������������������U����E�E��   �� �U��
%�  ��f�E��M����   uG3ҋEf��   �� �U��
��u�   k� �E����u	�E�   ��E�   f�E��j�h�U����E�P������f�E��M���>�   �� �E��������� ?  �   �� �E�f��M���~�Uf�
�����
3��Mf�3���]�����������������������������������������������������������U���V�   k��U�
% �  f�E��   f�M��   k��M����U��   k��Uf�E�f�
�M��u<�   ��E���u*�   �� �E���u�   k� �M����y  ��E���f�E��   k��E���un�   ��   k��E�uf�f��   �� �   ��U�uf�f�
�   k� �   �� �M�uf�f��   k� 3ҋEf��t����f�M�f��f�M��   k��M�����   �   k��U�
��   ��U�
����   k��Uf�
�   ���M���   �� �M���й   ��Ef��   �� �U�
��   k� �M���¹   �� �Uf�
�   k� �Uf�
f��   k� �Mf������f�U�f��f�U��   k��U�
�� ��   �   k� �E����   �� �E���ʸ   k� �Ef��   �� �U�
���   ��U�
����   �� �Mf��   ��E����   k��U���Ⱥ   ��Ef��   k��Ef�f��   k��Uf������   k��U�
���   k��Mf��   k��M��U���   k��Mf�f�E�^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�E��   k��E�����  ��f�M��U����  ug�   k��U��
��uA�   ��U��
��u/�   �� �U��
��u�   k� �E����u	�E�   ��E�   f�E��  �V�   k��M�������u?�   ���M����u-�   �� �M����u�   k� �U��
��u3��  �M��3  +��E+�f�U��M���3��  �  �U���5|b�   k��U��
% �  �   k��M�f��   ��3��M�f��   �� 3��M�f��   k� 3ɋU�f�����  �  �E���f�E\�f�M�f�U�f��f�U��E���|��U��J�M�#�f�M��U���|��M��U��B3��M���|��M�f�Q�U��U��}�t`�}�t0�}�t�|�   ���M���E��f�E��   ��3ҋE�f��   �� �U��
�M��f�M��   �� 3��M�f��   k� �M���E��f�E��   k� 3��M�f��U���t	�E�������E�    f�E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�E��   k��E�����  ��f�M��U����  ul3��Mf��   k��M����uA�   ���M����u/�   �� �M����u�   k� �U��
��u	�E�   ��E�   f�E��l�j�M����U�R�������f�E��E���@�   k��E����������?  �   k��U�f��E�-�  �Mf������
3ҋEf�3���]�����������������������������������������������������������������������������������U���EP�MQ�%�����]�����������U��EP�MQ�� ����]������������U��SV��څ�t��t�U��tW�̋�����F�^�2_^[]� ��������������U��QS�ډM�VW��tM3�93~G3����    �K�E��9�|�����u�D9U��<����t�t9�EP�������F��;3|Ëu3��ƅ�t`�@G��u���tT�>����u�~����u�~����u	�~����t�EWVP�y������F�|0�����t�EWVP�^������vO��u�_^[��]� ���������������������������������������������������������������U��QS�ډM�V3�93~AW3��K�E��9�|�����u�D9U��<����t�t9�EP�������F��;3|�_^[��]�������������������������u�U��� PRSVW�Ej P�������_^[ZX��]�����������̀=�� uj jj j j �������P�������������������������������jjj j j �b�������������������U����P�]����������������U��Q���P��E��}� t�U�j������jj ������^�����]����������������������U��Q�E�    ���P��E��MQ�����E���]�����������������U��Qh�   h��jjj �������E��E�P�����������}� u�   ��U��    3���]���������������������������U��j�hȒh�Ld�    P���SVW���1E�3�P�E�d�    �E�    �����E�    �EP�T   ���E��E������   �����ËE�M�d�    Y_^[��]��������������������������������������U������P��E����Q��E��U�;U�r�E�+E�����s3���   j�M�Q��������E�U�+U���9U���   �}�   s�E�E���E�   �M�M�M��U�;U�r"j}h��j�E�P�M�Q��������E�}� u:�U���U��E�;E�r%h�   h��j�M�Q�U�R��������E�}� u3��Q�E�+E����M���U��E�E��M�Q�����UR��M���U����U��E�P�����E��]����������������������������������������������������������������������������������U��Q�EP�$�������u	�E�������E�    �E���]����������������������U��� ���j��������EP��������=�� u
j�������h	 ��P�����]���������������������������U���$  j������t�   �)�������������5���=��f���f���f���f���f�%��f�-�������E ����E����E�����������  ���������	 ����   ���   �   k� ǂ��   �   k� ����T��   �� ����L�hȸ������]������������������������������������������������������������������������������U��j�,���]�����U���  j�V�����t�M�)�������������5���=��f���f���f���f���f�%��f�-�������E ����E����E������������������	 ����   ���   �   k� �E����hȸ�Q�����]���������������������������������������������������������������U���   j�F�����t�M�)�������������5���=��f���f���f���f���f�%��f�-�������E ����E����E������������������	 ����   �} v�} u�E    �}v	�M���M�U������   k� �U�����E�    �	�E����E��M�;Ms�U��E��M��������hȸ�������]����������������������������������������������������������������������������U��EP�MQ�UR�EP�MQ�I�����]����������������U��EP�MQ�UR�EP�MQ����]�������������������U���0  ���3ŉE��}�t�EP�J�����ǅ����    jLj ������Q��������������������0���������ǅ����    ǅ����    ������������������������������������f������f������f������f������f������f�������������ǅ0���  �M�������U�������E�H��������U�������E�������M������� ������������R�.����������������� u������ u�}�t�EP�$������M�3�������]����������������������������������������������������������������������������������������U��Q�E�    �x��E��M�Q��E��E���]����������U��E�x�]����U��Q�x��E��M�Q��E��}� t�UR�EP�MQ�UR�EP�U�����MQ�UR�EP�MQ�UR�5�����]�������������������������U��j������t�   �)jh �j�u�����h ��a�����]����������������������������U��Q�E�    �x��E��M�Q��E��UR��E�E�x��E���]���������������������U��j���E�$���E�$�D   ��]����������������U��j���E�$���E�$�   ��]����������������U���8Vh��  h?  �������E��E%�  =�  t�M���  ���  ��   �U���  ���  u�E����u(�} u"�M���  ���  uE�U����u�} t5�E�P�E�E���$���E�$���E�$�MQj�U�����$�b  �U���  ���  t�E%�  =�  u'�M�Q���E�$���E�$�UR�2������  h��  �E�P�������p���  ���]����Au�E���]���]����Au�E���]�E�]����z�E�]���E�]��E��]��E���������Dzh��  �M�Q�*��������  �E�u��]�E�u��]�E�M�E�M���]ЍU�R���E��$�0�  �$�a�����E�P���E��$�]��I�����M��]�u�u����E��$���������u��}�   ~P�M���   Q���E��$�������]�U�R���E��$���E�$���E�$�EPj讶����$�   �}����}M�M���   Q���E��$��������]�U�R���E��$���E�$���E�$�EPj�U�����$�e�M�Q���E��$�~������]�U��� th��  �E�P��������E��/�-�M�Q���E��$���E�$���E�$�URj������$^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�EP�x�����]��������������WV�t$�L$�|$�����;�v;��h  �%D�s��  ���   ��  ��3Ʃ   u�%ܺ��  �%D� ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf����s����   u������r*��$�s��Ǻ   ��r����$�,r�$�(s��$��r�<rhr�r#ъ��F�G�F���G������r���$�s�I #ъ��F���G������r���$�s�#ъ���������r���$�s�I s�r�r�r�r�r�r�r�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�s��(s0s<sPs�D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$��t�����$�dt�I �Ǻ   ��r��+��$��s�$��t��s�st�F#шG��������r�����$��t�I �F#шG�F���G������r�����$��t��F#шG�F�G�F���G�������V�������$��t�I htptxt�t�t�t�t�t�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��t���t�t�t�t�D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} u3��  �} t	�E�   ��E�    �E��E��}� u#hԸhpjj j7h�j葭������u̃}� u0������    j j7h�hX�hԸ�4������   �6  �} t�U;U�  �EPj �MQ�A������} t	�E�   ��E�    �U�U��}� u#hp�hpjj j=h�j��������u̃}� u0�G����    j j=h�hX�hp��������   �   �M;Mr	�E�   ��E�    �U�U�}� u#h��hpjj j>h�j�u�������u̃}� u-������ "   j j>h�hX�h���������"   ��   ��MQ�UR�EP�m�����3���]������������������������������������������������������������������������������������������������������������������������̋T$�L$��t�D$�%D�s�L$W�|$��]�T$���   |�%ܺ�,���W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$������������������������������������������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+���������������������������������������WV�t$�L$�|$�����;�v;��h  �%D�s��  ���   ��  ��3Ʃ   u�%ܺ��  �%D� ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf�����~����   u������r*��$��~��Ǻ   ��r����$��}�$��~��$�<~��}�}~#ъ��F�G�F���G������r���$��~�I #ъ��F���G������r���$��~�#ъ���������r���$��~�I �~�~�~|~t~l~d~\~�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��~���~�~�~�~�D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$�D������$���I �Ǻ   ��r��+��$�H�$�D��X|��F#шG��������r�����$�D��I �F#шG�F���G������r�����$�D���F#шG�F�G�F���G�������V�������$�D��I � ���� �(�;��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�D���T�\�l����D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M��EP�M��؝���M����E���]� �����������U��Q�M��EP�M��R����M����E���]� �����������U��Q�M��EP�M��?����M����E���]� �����������U��Q�M��EP�M������M����E���]� �����������U��Q�M��EP�M�������M�����E���]� �����������U��Q�M��EP�M�芴���M�����E���]� �����������U��Q�M��E�� Ĺ�M��A    �U��B �E�Q�M������E���]� ������������������������U��Q�M��E�� Ĺ�M��U��A�M��A �E���]� ���������������������U��Q�M��E�� Ĺ�M��A    �U��B �EP�M������E���]� ��������������������������U��Q�M��E�� Ĺ�M��A    �U��B �E���]�������������������������U��Q�M��E�� ��M��#�����]���������������������U��Q�M��E�� ��M�������]���������������������U��Q�M��E�� ���M�������]���������������������U��Q�M��E�� Ĺ�M��������]���������������������U��Q�M��E�;Et0�M������M�Q��t�E�HQ�M��0�����U��E�H�J�E���]� ������������������������U��Q�M��M������E��t�M�Q�@������E���]� ��������������������U��Q�M��M��V����E��t�M�Q� ������E���]� ��������������������U��Q�M��M�茪���E��t�M�Q��������E���]� ��������������������U��Q�M��M��k����E��t�M�Q�������E���]� ��������������������U����M��} tK�EP����������E��M�Q� ������U��B�E��x t�MQ�U�R�E��HQ�?������U��B��]� ��������������������������������U��Q�M��E��H��t�U��BP�������M��A    �U��B ��]���������������������������U����M��E��x t�M��Q�U���E�й�E���]����������������������U����E������} t	�E�   ��E�    �E�E��}� u#h��hpjj jYh@�j藜������u̃}� u.������    j jYh@�hԺh���:���������   �U�U��E��H��   ta�U�R��������E��E�P�p������M�Q������P�D�������}	�E������$�U��z tj�E��HQ蘪�����U��B    �E��@    �E���]���������������������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E������} t	�E�   ��E�    �E�E��}� u#h�hpjj j.h@�j��������u̃}� u+�r����    j j.h@�h��h������������W�U�B��@t�M�A    �=�UR�������E�    �EP荸�����E��E������   ��MQ�������ËE܋M�d�    Y_^[��]���������������������������������������������������������������������������U��Q�} uj �_  ���S�EP��������t����>�M�Q�� @  t.�EP�V�����P��������t	�E�������E�    �E��3���]������������������������������������U����E�    �E�E��M��Q����u|�E��H��  tn�U��E��
+H�M��}� ~Z�U�R�E��HQ�U�R������P�Ͼ����;E�u�E��H��   t�U��B����M��A��U��B�� �M��A�E������U��E��H�
�U��B    �E��]��������������������������������������������������������U��j��   ��]������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} uj �   ���@�EP�������E�    �MQ�i������E��E������   ��UR�D�����ËE�M�d�    Y_^[��]������������������������������������������������������U��j�h(�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    j�u������E�    �E�    �	�E���E�M�;���   �U䡜�<� ��   �M�����H��   ��   �U䡜��Q�U�R躳�����E�   �E�����B%�   te�}u%�M����P���������t	�M����M��:�} u4�U䡜���Q��t!�E����R�֨�������u�E������E�    �   ��E����R�E�P�<������������E������   �j������Ã}u�E����E܋M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������U����E�H���M��U�E��B�}� |�M��%�   �E��M����E���MQ�������E��E���]���������������������������U��j�hX�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E܉E؃}� u#h�hpjj j)h��j�͔������u̃}� u.�"����    j j)h��hX�h��p���������  �UR��������E�    �E�EԋMԋQ��@��   �E�P��������E�}��t!�}��t�M����U�����P��U���E���EЊH$�����х�uA�}��t!�}��t�E����M�����P��M���E���ŮB$�� ���ȅ�t	�E�    ��E�   �UȉUă}� u#hh�hpjj j-h��j裓������u̃}� u-������    j j-h��hX�hh��F������E������}� uP�M�Q���U��E�M��H�}� | �U�����   �M��U����M���UR��������E��E��E��E������   ��MQ�0�����ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hx�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E܉E؃}� u#h�hpjj jCh��j�͑������u̃}� u.�"����    j jCh��h��h��p���������  �UR��������E�    �E�EԋMԋQ��@��   �E�P��������E�}��t!�}��t�M����U�����P��U���E���EЊH$�����х�uA�}��t!�}��t�E����M�����P��M���E���ŮB$�� ���ȅ�t	�E�    ��E�   �UȉUă}� u#hh�hpjj jGh��j裐������u̃}� u-������    j jGh��h��hh��F������E������}� uP�M�Q���U��E�M��H�}� | �U�����   �M��U����M���UR��������E��E��E��E������   ��MQ�0�����ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u#h�hpjj j-h��j���������u̃}� u.�S����    j j-h��h�h�����������   �} t	�E�   ��E�    �U�U��}� u#h �hpjj j.h��j腎������u̃}� u+������    j j.h��h�h ��(���������3�MQ��������M��Q�U�U�E�M�#Q���t3��������]�������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E܉E؃}� u#h��hpjj j,hH�j�M�������u̃}� u.�����    j j,hH�h��h�������������  �UR�S������E�    �E�EԋMԋQ��@��   �E�P�G������E�}��t!�}��t�M����U�����P��U���E���EЊH$�����х�uA�}��t!�}��t�E����M�����P��M���E���ŮB$�� ���ȅ�t	�E�    ��E�   �UȉUă}� u#hh�hpjj j0hH�j�#�������u̃}� u-�x����    j j0hH�h��hh���������E������}� uZ�M�Q���U��E�M��H�}� |&�U��M��U���   �U��E����U�
��EP�MQ��������E��U��U��E������   ��EP������ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E܉E؃}� u#h��hpjj jGhH�j�=�������u̃}� u.�����    j jGhH�h��h�������������  �UR�C������E�    �E�EԋMԋQ��@��   �E�P�7������E�}��t!�}��t�M����U�����P��U���E���EЊH$�����х�uA�}��t!�}��t�E����M�����P��M���E���ŮB$�� ���ȅ�t	�E�    ��E�   �UȉUă}� u#hh�hpjj jKhH�j��������u̃}� u-�h����    j jKhH�h��hh��������E������}� uZ�M�Q���U��E�M��H�}� |&�U��M��U���   �U��E����U�
��EP�MQ��������E��U��U��E������   ��EP������ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u#h�hpjj j*hȽj�^�������u̃}� u.�����    j j*hȽh,�h�����������   �} t	�E�   ��E�    �U�U��}� u#h �hpjj j+hȽj��������u̃}� u+�:����    j j+hȽh,�h �����������j �M�QR�P�MQ舔������]��������������������������������������������������������������������������������U��j�hؓh�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h�hpjj j;h@�j�ͅ������u̃}� u.�"����    j j;h@�h��h��p����������   �} t�}t�}t	�E�    ��E�   �U܉U؃}� u#h��hpjj j<h@�j�H�������u̃}� u+�����    j j<h@�h��h�������������L�MQ�Q������E�    �UR�EP�MQ�UR�f������E��E������   ��EP�������ËEԋM�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������U����} u#hl�hpjj jch@�j��������u̋M�M��U��B%�   t�} t�}t�}t�P����    �����   �M��Q���E��P�}u�M�Q腪����EU�E�U�E    �U�R�&������E��H��   t�U��B����M��A�.�U��B��t#�M��Q��t�E��H��   u
�U��B   �EP�MQ�UR�E�P蟶����P�?������E��U�M�#M���u	�E�������E�    �E���]������������������������������������������������������������������������������������U���H�} t�} u3���  �} t	�E�   ��E�    �E�E��}� u#h�hpjj jqh��j�[�������u̃}� u-�����    j jqh��h��h��������3��t  �} t	�E�   ��E�    �U܉U؃}� u#h�hpjj jrh��j��������u̃}� u-�8����    j jrh��h��h�������3���  ���3��u9Ew	�E�   ��E�    �MԉMЃ}� u#hD�hpjj jsh��j�d�������u̃}� u-�����    j jsh��h��hD�������3��}  �E�E�M�M�M��U��U��E�H��  t�U�B�E���E�   �}� �:  �M�Q��  ��   �E�x ��   �M�y }N�U�z }&h��hpjj h�   h��j蚀������u̋M�Q�� �E�P�E�+E�3��u��  �M�U�;Qs�E��E��	�M�Q�ŰẺE��M�Q�U�R�E�Q艉�����U�+U��U��E�H+M��U�J�E�M��U�
�E�E��E��T  �M�;M���   �U�B%  t �MQ�o�������t�E�+E�3��u�#  �}� t�E�3��u�E�+E���M��MȋUȉU��E�P�M�Q�UR������P�������E�}��u�E�H�� �U�J�E�+E�3��u�   �E�;E�v�M��M���U�UċEĉE��M�+M��M��U�U��U�E�;E�s�M�Q�� �E�P�E�+E�3��u�h�^�M���U��EP�M�Q�M��������u�E�+E�3��u�;�U���U�E����E��M�y ~�U�B�E���E�   �M��M������E��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t�} u3���   �} t	�E�   ��E�    �E�E��}� u#h�hpjj jMh��j�}������u̃}� u*�o����    j jMh��h�h�轻����3��L�UR�$������E�    �EP�MQ�UR�EP�/������E��E������   ��MQ�ҹ����ËE܋M�d�    Y_^[��]������������������������������������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E��E܃}� u#h��hpjj j6h`�j�{������u̃}� u.�����    j j6h`�h��h���`���������/  �}t�} t�}@t	�E�    ��E�   �U؉Uԃ}� u#h��hpjj j<h`�j�8{������u̃}� u.�����    j j<h`�h��h���۹��������  �} t
�}@��   �}r�}���w	�E�   ��E�    �MЉM̃}� u#h`�hpjj j@h`�j�z������u̃}� u.������    j j@h`�h��h`��I���������  �E����E�M�M�U�R蝰�����E�    �E�P�Ƚ�����M�Q�t������U�B%�����M�A�U��t!�E�H���U�J�E���E�E   �b�} uJjxh��j�MQ��u�����E�} u�|����|��E������J�E�H��  �U�J��E�H��   �U�J�E�M�H�U�E�B�M�U��E��@    �E������   ��M�Q莶����ËEȋM�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���$�E�E�M�Q��@��   �E�P�ī�����E��}��t!�}��t�M����U������P��U���E���E��H$�����х�uA�}��t!�}��t�E����M������P��M���E���U�B$�� ���ȅ�t	�E�    ��E�   �U�U�}� u#hh�hpjj j#hX�j�w������u̃}� u.������    j j#hX�h��hh��C���������  �M�M��}�t$�U��B��u!�M��Q��   t�E��H��t�����   �U��z u�E�P�հ�����M��U��;Bu�M��y t����   �U�����M���U��B��@t5�M�����U��E��M���U���M;�t�U�����M������R��U�����E܋M��U܉�E܊M��U��B���M��A�U��B���M��A�U��B���M��A�E%�   ��]��������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h8�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h�hpjj j/h��j�Mu������u̃}� u+袻���    j j/h��hH�h�����������D�UR�V������E�    �EP�MQ�J������E��E������   ��UR������ËE܋M�d�    Y_^[��]������������������������������������������������������������������������������U��Q�=� u��   ��=�}
��   h�   h��jj��P詌�������=� u<��   h�   h��jj��Q�t��������=� u�   �3�E�    �	�U����U��}�}�E���`��M�������3���]��������������������������������������������������������U�����������t��v��j��Q���������    ]����������������������������U��`�]�������U��}`�r?�    k���`�9Mw,�U��`�����R��s�����E�H�� �  �U�J��E�� P� ]�����������������������U��}}#�E��P�s�����M�Q�� �  �E�P��M�� Q� ]����������������������U��}`�r>�    k���`�9Mw+�U�B%����M�A�U��`�����R�^�������E�� P�]������������������������U��}}#�E�H������U�J�E��P��������M�� Q�]����������������������U����E�E��M�Q�UR�EP�MQ�UR�EP�MQ�������E��E�    �E���]��������������������������������U����E�E��M�Q�UR�EP�MQ�UR�EP�MQ�w�����E��E�    �E���]��������������������������������U��E P�MQ�UR�EP�MQ�UR�EP虫����]������������������������U��j�hX�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t�}t	�E�    ��E�   �E܉E؃}� u#h��hpjj jth�j�p������u̃}� u.�l����    j jth�hp�h��躮��������  �} t	�E�   ��E�    �UԉUЃ}� u#h��hpjj juh�j�o������u̃}� u.�����    j juh�hp�h���A���������  j�Tp�����E�    �D��M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���M̋U�ẺB�M̉M��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H�D�j�U�R�W}�����<3�u&h��hpjj h�   h�j�n������u��E������ߴ���    ��   �}� tu�U�B���EȋM�UȉQ�EȉE��M�;D�tM�U�z t�E�H�U���M��E�H�J�U��    �E�D��H�D��E��M�D��h�   h<�jj��i�����E�}� u�E������.����    �L�U��    �E�D��H�=D� t�D��E��M��A   �E�   �U�E�B�M�D��E������   �j详����ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��\"  �R������3ŉE�ǅ����    ǅ����    ǅ����    �} u
�   �S  ������P�MQj�,��u
ǅ����    �   i�  ������������
  s������3ɋ�����f������h  ������P������Q�(��u8j h_  h�hl�h��h�h  ������R�Ͳ����P�`v����������������������Q��������@vo������R�������������TA�������j hh  h�hl�hX�j�`�P������������+����  +���P������Q�w����P��u�����} t*�UR葔������@v�EP耔�����M�TA��������&���� �����������     �}uǅ����h��
ǅ����p��   k� �E���t�U�������
ǅ����p��   k� �U�
��t�}uǅ����|��
ǅ����p��   k� �E���tǅ�������
ǅ����p��} t�U�������
ǅ����p��} tǅ�������
ǅ����p��} t�E�������
ǅ����p��} tǅ�������
ǅ����p������� t�������������'�} t�U�������
ǅ����p������������������� tǅ����t��
ǅ����p��} tǅ�������
ǅ����p�������Q������R������P������Q������R������P������Q������R������P������Q������R������P�M���Rh��h�  h   ������P�{�����D������������ }*j h  h�hl�h��j"j�����Q��e���� �ծ��������������� }8j h�  h�hl�h��h��h   ������P�o�����P�s����h  h��������Q觇����������������uj��u����j��i��������u�   �3��M�3�蛆����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��} u��EP�MQ�UR�EP�MQ�Ť��]�����������U��} t�E;Et�M;Mt�E��U$R�E P�MQ�UR�EP肤���E]���������������������U��Q�M��E��@ �} ��   �D����M��A�U��B�M��Pl��E��H�U��Ah�B�M��;4�t�E��H�Qp# �u
贠���M���U��B;|�t�M��Q�Bp# �u�أ���M��A�U��B�Hp��u�U��B�Hp���U��B�Hp�M��A��U��J�U���J�E���]� ���������������������������������������������������������U��Q�M��E��H��t�U��B�Hp����U��B�Hp��]����������������������U��Q�M��E���]�������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j�le�����E�    h��hDtj j j j �d������u̃} t�M��U࡜��E���M��U�}� �0  �E�;E��$  �M�Q����  ��t)�E�H����  t�U�B%��  ��u�l���u��  �U�z tyj j�E�HQ���������tj�U�BP��  ����t$�M�QRh��j j j j ��c������u��)�M�QR�E�HQh��j j j j �c������u̋E�HQh��j j j j �c������u̋E�H����  ����   �U�BP�M�Q������  R�E�� Ph��j j j j �Nc���� ��u̃=�� t3�U�BP�M�� Q��  ����u�U�BP�M�� Q�������U�R�EP�7  ���   �M�yu;�U�BP�M�� Qh0�j j j j ��b������u̋E�P�MQ�A7  ���Y�U�B%��  ��uI�M�QR�E�H������  Q�U�� Rh`�j j j j �pb���� ��u̋M�Q�UR��6  �������E������   �j�,������h��hDtj j j j �"b������u̋M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hؕh�Ld�    P���SVW���1E�3�P�E�d�    �e��E�    3��E��E��E��E��EĉEȉẺEЍM�Q�4�U��U؃} ��   �} u
�   �   �E�E��M�U��D
��E܋M�;M�s	�   �v�r�E�    �U���E�M؃���#M��M��U؃���#U܉U܋E�;E�t�M�M؉M��U���E����E������#�   Ëe��E�   �E������E��	�E�����3��M�d�    Y_^[��]�����������������������������������������������������������������������������������������U����E�E��M���M�}� t'�U��E��M�M�U���U�E�;E�t3���ĸ   ��]����������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�   �l���u
�   ��  j�_�����E�    �Ї���Eԃ}����   �}����   �MԉM܋U܃��U܃}���   �E��$���h �hDtj j j j �^������u��   h,�hDtj j j j �^������u��dhX�hDtj j j j �k^������u��Bh��hDtj j j j �I^������u�� h��hDtj j j j �'^������u��E�    ��  ����E���M��U�}� ��  �E�   �E�H����  ��t#�U�zt�E�H����  ��t	�U�zu�E�H����  ��P��U���E���j�t�P�M��Q���������uz�U�z t=�E�HQ�U�BP�M�� Q�U�BP�M�Qh��j j j j �D]����(��u��-�E�� P�M�QR�E�Ph��j j j j �]���� ��u��E�    j�t�R�E�H�U�D
 P�$�������uz�M�y t=�U�BP�M�QR�E�� P�M�QR�E�Ph8�j j j j �\����(��u��-�U�� R�E�HQ�U�Rh �j j j j �w\���� ��u��E�    �M�y ��   �U�BP�v�Q�U�� R�{�������ud�E�x t2�M�QR�E�HQ�U�� Rh��j j j j �\���� ��u��"�M�� Qh��j j j j ��[������u��E�    �}� uz�E�x t=�M�QR�E�HQ�U�BP�M�� Q�U�RhH�j j j j �[����(��u��-�M�QR�E�� P�M�Qh��j j j j �d[���� ��u��E�    �G����E������   �j�)�����ËEЋM�d�    Y_^[��]Ð����`�;���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h8�h�Ld�    P���SVW���1E�3�P�E�d�    �} t	�E�   ��E�    �E��E܃}� u&h��hpjj h�  h��j�!Y������u̃}� u+�v����    j h�  h��h��h����������s�l���u�fj��Y�����E�    ����E���M��U�}� t$�E�H����  ��u�UR�E�� P�U�����E������   �j�ˑ����ËM�d�    Y_^[��]�����������������������������������������������������������������������������������U���8���3ŉE��E�P��������   ���|� u'�   �� �|� u�l���t?�   ��|� t1h��hDtj j j j �X������u�j �H������   �3��M�3��Nv����]����������������������������������������������U��h�]�������U�졀�]�������U�졈�]�������U��j�hX�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�     �} t	�M�    �} t	�U�    �EP�3������u3���   j�W�����E�    �M�� �M�U�B%��  ��t"�M�yt�U�B%��  ��t	�M�yukj�UR�EP�J�������tU�M�Q;UuJ�E�H;p�<�} t�U�E�H�
�} t�U�E�H�
�} t�U�E�H�
�E�   ��E�    �E������   �j������ËE��M�d�    Y_^[��]���������������������������������������������������������������������������������������������������U��} u3��1j j �E�� P�:�������u3���M�� Qj ���R�0]�����������������U��Q�} t	�E�   ��E�    �E���]����������������U��j�hx�h�Ld�    P���SVW���1E�3�P�E�d�    �} t	�E�   ��E�    �E܉E؃}� u&h�hpjj h�  h��j�aT������u̃}� u.趚���    j h�  h��h@�h��������m  j�U�����E�    �U�����E�    �	�M����M��}�}�U��E�D�    �M��U�D�    �ӡ���E���M��U�}� ��   �E�H����  |f�U�B%��  ��}V�M�Q����  �E�L����U�B%��  �U�L��E�H����  �U�D��M�A�U�J����  �U�D��W�E�x t/�M�QR�E�HQ�U�Rhl�j j j j �zS���� ��u���M�Qh��j j j j �YS������u������E����H,�U����B0�E������   �j������ËM�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������U��� V�E�    �} t	�E�   ��E�    �E��E�}� u&h�hpjj h�  h��j��Q������u̃}� u0�����    j h�  h��h��h��c�����3���  �} t	�E�   ��E�    �U��U�}� u&h�hpjj h�  h��j�EQ������u̃}� u0蚗���    j h�  h��h��h�������3��E  �} t	�E�   ��E�    �M�M�}� u&h4�hpjj h�  h��j��P������u̃}� u0�����    j h�  h��h��h4��g�����3���   �E�    �	�E����E��}�}�M��U�E��u�L�+L��U��E�L��M��U�E��u�L�+L��U��E�L��M��U�|� u�E��M�|� t$�}� t�}�u�}�u�l���t�E�   �r����E�M�P,+Q,�E�P,�M�U�A0+B0�M�A0�U�    �E�^��]�������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    �E�P�M���X���M��%���P�MQ�E������M��i����]�����������������������U����} t	�E�   ��E�    �E��E�}� u&h�hpjj h
  h��j�N������u̃}� u.������    j h
  h��h��h��+������   �E�    �	�U����U��}�}>�E���P�Q�U��E�L�Q�U��E�L�Qh�j j j j �gN���� ��u�볋E�H,Qh,�j j j j �CN������u̋E�H0QhT�j j j j �!N������u̋�]���������������������������������������������������������������������������������U��Q�EP��u������u�����M�� �M��U��B��]���������������������U��Q�h��E��M�h��E���]���������������������U��Q�d��E��M�d��E���]���������������������U��Q����E��E���]��������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    j�cM�����E�    �EP��t������tj�M�� �M�U�B%��  ��tH�M�yt?�U�B%��  ��t/�M�yt&h`�hpjj h?  h��j��K������u̋E�M�H�E������   �j�#�����ËM�d�    Y_^[��]�����������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �l��E܃}�t�M����  ���t	�E�    ��E�   �U�U��}� u&h��hpjj hw  h��j��J������u̃}� u0�P����    j hw  h��h��h��蛉�����l��sj�K�����E�    �l��M܃}�t7�U��t���   ��E��%��  ������    �M�l��E������   �j裃����ËE܋M�d�    Y_^[��]����������������������������������������������������������������������������������������U��Q�h��E��M�h��E���]���������������������U��Q����E��M����E���]���������������������U��EP�nc����]����������������U��Q�} u�   �E������E�j�t�Q�U��R���������t!�EPh�j j j j�vI������u��Lj�u�R�E���P��������u�MQh��j j j j�8I������u�j�E��Q�dW������]��������������������������������������������������������U��j j j �EP�MQ�I����]����������������������U��EP�MQj �UR�EP��H����]������������������U��EP�MQ�UR胔����]��������U���$�E�    �E�    �E�    �E�    �E�    �} t	�E�   ��E�    �E�E��}� u&hl�hpjj h  h��j�G������u̃}� u.�����    j h  h��h��hl��8���������w�E�    �U������U��E��Q��P�����E�U��E+�E�3�+M���M�}v�U�U���E�   �E���E�M�U�D
+E��E��M�+M�+M��M܋E܋�]���������������������������������������������������������������������������������U��j j �EP�MQ�UR�'G����]��������������������U���,�E��#Eu	�E�   ��E�    �M��M�}� u&h|�hpjj h@  h��j�F������u̃}� u0�k����    j h@  h��h��h|�趄����3��E  �} t�E;Er	�E�    ��E�   �M��M�}� u&h��hpjj hA  h��j�E������u̃}� u0�����    j hA  h��h��h���0�����3��   �}v�E�E���E�   �M���M3�+U���U܋E�M܍T�U��EE��E�M;M�v�n����    3��i�UR�EPj�M�Q��@�����E��}� u3��F�U�U�U�E��#�+U�UԋM�+M܃��M�j�u�R�E؃�P�k�����M؋U���Eԋ�]�������������������������������������������������������������������������������������������������������������������������������U��j j �EP�MQ�UR�EP躑����]����������������U���8�} u!�EP�MQ�UR�EP�MQ�jD������  �} u�UR�]����3��  �E������E�j�t�Q�U��R��������t1�EPh0�j j j j�C������u�趉���    3��_  j�u�R�E���P���������u�MQh��j j j j�qC������u̋E��#Eu	�E�   ��E�    �M��M�}� u&h|�hpjj h�  h��j��B������u̃}� u0�����    j h�  h��h��h|��`�����3��  �} t�E;Er	�E�    ��E�   �M�M�}� u&h��hpjj h�  h��j�:B������u̃}� u0菈���    j h�  h��h��h���ڀ����3��  �E��Q�K�����U��M+
+��Ẽ}v�U�U���E�   �E����E3�+M���MԋU�EԍL�M؋UU؉U܋E;E�v������    3��   �MQ�URj�E�P�=�����E��}� u3��   �M�M�M�U��#�+M�M�E�+Eԃ��E�j�u�Q�UЃ�R�9h�����EЋM���U�;Uv�E�E���M̉MȋU�R�EP�M�Q�CJ����j�U��P�O�����E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j j �EP�MQ�UR�EP�MQ��G����]������������U����E�    �E�    �E�    �} v�����3��u;Es�����    3��s�E�E�E��} t�MQ�UR�EP�������E��M Q�UR�EP�MQ�U�R�EP�#������E�}� t �M�;M�s�U�+U�Rj �E�E�P�Df�����E��]�����������������������������������������������������������U��j j j �EP�MQ�UR蜌����]������������������U��EP�MQj �UR�EP�MQ�h�����]��������������U��j j j �EP�MQ�UR�EP�BF����]��������������U��EP�MQj �UR�EP�MQ�UR�F����]����������U����E�    �E�P�MQ�UR�EP�MQ�UR�[f�����E��}� u�}� t�X�����t
�O����M���E���]���������������������������U��Q�} v�����3��u;Es�����    3��K�E�E�E�MQ�UR�EP�MQ���R�EP��  ���E��}� t�MQj �U�R�cd�����E���]������������������������������������������U��Qj j j�EP�MQ�XR�����E��E���]�������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E��E܃}� u&h��hpjj h�  h��j�z<������u̃}� u-�ς���    j h�  h��h��h���{����3��c�}�v蜂���    3��Nj�=�����E�    j �UR�EP�MQ�UR�EP��  ���E��E������   �j�5u����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������U��j�h��h�Ld�    P��SVW���1E�3�P�E�d�    j�C<�����E�    �EP�MQ�Zm�����E������   �j�mt����ËM�d�    Y_^[��]�������������������������������������U��Q�=�� vZ�����9��u;��Y����u&h��hpjj h  h��j�:������u����    ����������} u�  �}uOj�u�P�M�����Q���������t/�URh��j j j j�:������u�荀���    �5  �=h� tDj j j �MQj �URj�h�����u%h@�hDtj j j j �>:������u���  �MQ�Jb������u&hh�hpjj h*  h��j�9������u̋E�� �E��M��Q����  ��tI�E��xt@�M��Q����  ��t/�E��xt&h`�hpjj h0  h��j�<9������u̋l����m  j�t�P�M���Q����������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��P�Ph��j j j j�9����(��u��<�U��� R�E��HQ�U��B%��  ��P�Qh��j j j j��8���� ��u�j�t�P�M��Q�E��L Q�����������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��P�Ph8�j j j j�b8����(��u��<�U��� R�E��HQ�U��B%��  ��P�Qh �j j j j�$8���� ��u̋E��xuj�M��y����u	�U��z t&h��hpjj hi  h��j�|7������u̋M��Q��$R�v�P�M�Q�h^�����U�R��o�����`  �E��xu�}u�E   �M��Q;Ut&h4�hpjj hw  h��j�7������u̋M����+Q����l�����   �M��9 t�U���M��Q�P�;���;E�t&h|�hpjj h�  h��j�6������u̋U��B����M��y t�U��B�M����:���;E�t&h��hpjj h�  h��j�K6������u̋U������M��Q��$R�v�P�M�Q�-]�����U�R�n�����(�E��@    �M��QR�v�P�M��� Q��\������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�EP�f����]��������������U��j j j�EP�\i����]����������U����E�    �E�P�MQ�UR�EP�MQ�J   ���E��}� u�}� t�z����t
�z���U���E���]�������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    j�4�����E�    �=�� vZ�����9��u;�R����u&h��hpjj h  h��j�b3������u����    ����������p��E��=d��t�M�;d�u̃=h� tu�UR�EP�M�Q�UR�EPj j�h�����uP�} t%�MQ�URh�j j j j �73������u�� hX�hDtj j j j �3������u��D  �U����  ��t�l���u�E�   �}�v3�MQh��j j j j��2������u̃} t	�E�    ��  �M����  ��t:�}t4�U����  ��t&�}t h��hDtj j j j�p2������u̋M��$�MԋU�R�#P�����E�}� u�} t	�E�    �r  �p����p��}� tI�U��    �E��@    �M��A    �U��B�����E�M�H�U��B   �E��@    �   ���+��;Mv���U����
����������E������;��v�������=�� t����M�H�	�U����E�����U��B    �E�M�H�U�E�B�M�U�Q�E�M�H�U�E��B�M���j�t�R�E��P�W����j�t�Q�U�E�L Q�W�����UR�w�P�M�� Q�{W�����U�� �U��E������   �j�i����ËE؋M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�EP�MQ�UR���P�MQ�j�����E��E���]���������������������U��j�EP�[����]��������������U��j�hؔh�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E��E܃}� u&h��hpjj h�  h��j�j.������u̃}� u1�t���    j h�  h��h��h���
m��������G  �=�� v[�����9��u;�FM����u&h��hpjj h�  h��j��-������u����    ���������j�.�����E�    �UR�3V������u&hh�hpjj h�  h��j�-������u̋M�� �M�U�B%��  ��tH�M�yt?�U�B%��  ��t/�M�yt&h`�hpjj h�  h��j�'-������u̋E�xu�}u�E   �M�Q�U��E������   �j�=f����ËE؋M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������U��j j j�EP�MQ�&g����]����������������������U����E�    �E�P�MQ�UR�EP�MQ�UR�F   ���E��}� u�}� t�8r����t
�/r���M���E���]���������������������������U��Q�EP�MQ�UR�EP�MQ�������E��}� t�E��?�} u�} t	�U�   �E��%�EP��c������u�} t	�M�   3��뗋�]��������������������������������U���x���3ŉE��EP�M���4���E�    �	�M����M��U�z}�E�H�M���E�   �U�;U���   �EE��H �M��M���w����t0�M���w����zt~ �M��w��PhW  �E�P�>�����E��hW  �M�Q�M��w��P�2&�����E��}� t	�U��U���E�    �E��M��L��p����U��p���     �E�Ph\�kM��1   +�RkE��L�Q�+d������}*j h	  h��hd�h��j"j�?p���R�0'���� �/p���M��������U��U��}�s��h���E��D� �M�Q�U�Rh��j j j j ��)������u̍M��C���M�3��9H����]�������������������������������������������������������������������������������������������������������������������������U��j�hx�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j�)�����E�    j�EP�MQ�UR�EP�MQ�}  ���E��E������   �j��a����ËE�M�d�    Y_^[��]������������������������������������������U��Qj j j�EP�MQ�UR��o�����E��E���]�������������������������U����E�    �E�    �E�    �} v�����3��u;Es�$n���    3��g�E�E�E��} t�MQ�41�����E��UR�EP�MQ�U�R�EP�x<�����E�}� t �M�;M�s�U�+U�Rj �E�E�P�`N�����E��]�������������������������������������������������������U����E�    �E��M��} u�UR�EP�MQ�U�R��"������  �} t�}� u�EP�MQ�e5����3��  �=�� v[�����9��u;��E����u&h��hpjj h�  h��j�u&������u����    ����������p��U�=d��t�E�;d�u̃=h� ty�MQ�UR�E�P�MQ�U�R�EPj�h�����uR�} t%�MQ�URh��j j j j �G&������u�� h,�hDtj j j j �%&������u�3��  �}��v`�} t)�UR�EP�M�QhX�j j j j��%���� ��u���E�Ph��j j j j��%������u���k���    3��A  �}th�U����  ��tZ�E%��  ��tM�} t%�MQ�URh��j j j j�n%������u�� h��hDtj j j j�L%������u��Qj�u�R�E�����P�d�������t1�MQh�j j j j�%������u��k���    3��  �EP�
M������u&hh�hpjj h  h��j�_$������u̋U�� �U�E�xu�E�   �}� t=�M�y����u	�U�z t&h��hpjj h#  h��j�$������u��d�M�Q����  ��u�E%��  ��u�E   �M���;Qs1�EPhh�j j j j�$������u��j���    3��  �} t%�U���$R�E�P�hr�����E��}� u3��c  �#�M���$Q�U�R�D�����E��}� u3��>  �p����p��}� u{�=���s;�M����+Q������+��;E�v���M�����
��������U����+B������M�������;��v
�������M��� �M�U��E�;Bv$�M��U�+QR�w�P�M��U�QR�I����j�t�P�M�M�Q�|I�����}� u�U��E�B�M��U�Q�E��M�H�U��E��B�} u4�} u�M�;M�t&h��hpjj h�  h��j�"������u̋E�;E�t�}� t�E���   �M��9 t�U���M��Q�P�;���;E�t&h �hpjj h�  h��j�!������u̋U��B����M��y t�U��B�M����:���;E�t&h\�hpjj h�  h��j�]!������u̋U������=�� t����U��Q��E�����M������E��@    �M�����E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;��u���RH�������������������U���,VW�   ����}��E�E��}� t:�M����t0�E��M��U����U��E��E�M��B�E��M�Q�U��H �ыU�U�E��E��}� t�M����t�E� @��E�P�M�Q�U�R�E�P�8_^��]� ��������������������������������������������������U��Q��E�H3M�J=��j �MQ�U�BP�M�QRj �EP�M�QR�EP�O^���� �E��E���]�����������������������U��QS��E�H3M��<���M�Q��ft�E�@$   �   �v�tj�M�QR�E�HQ�U�BPj �MQ�U�BP�MQ��]���� �U�z$ u�EP�MQ��]��j j j j j �U�Rh#  ������E��]�c�k ��   [��]������������������������������������������������������U����E�    �E�����M�3��E�U�U��E�E�M���M�d�    �E�E�d�    �UR�EP�MQ�l���E��E�d�    �E���]�������������������������������������XY�$�����������XY�$�����������XY�$�����������U���8S�}#  u��	�M��   ��   �E�    �E�p����M�3��EЋU�UԋE�E؋M�M܋U �U��E�    �E�    �E�    �e�m�d�    �EȍE�d�    �E�   �E�E��M�M��5N�����   �U��E�P�M�R�U����E�    �}� td�    ��]ȉd�    �	�E�d�    �E�[��]�����������������������������������������������������������������������U����MSVW�q�ދ}�A�E��u���x>�M���u�f���M�U�N��9L��U�}�U�;L��U�~���uO�u��څ�yȋM�EF�0�E�;Yw;�v�tf���M���_^[����]�����������������������������������������U��QS�E���E�d�    �d�    �E�]�m��c���[��]� ��������������U���SVWd�5    �u��E�^j �EP�M�Q�UR�<�E�H����U�Jd�=    �]��;d�    _^[��]� �����������������������U��MV�u��0L�����   �N�"L�����   ��^]�����������������������U��V��K���u;��   u��K���N^���   ]���K�����   �y t�A;�t�ȃy u�^]� e���F�A^]����������������������������U���K�����   ��t�M9t�@��u��   ]�3�]����������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ��X���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�X���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�@X���� �E�_^[�E���]���������������������U��E�HQ�   k� �M�T(Rj �E�HQ�����]� ����������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ����������������������������U��Q�M��E�� ���E���]� �������U��Q�M��E�� ���M�Q�[@������]�����������������U��Q�M��E���]� ����������������U����M��E���	P�M��	Q�uA������t	�E�    ��E�   �E���]� ��������������������U����M��E���	P�M��	Q�%A������t	�E�   ��E�    �E���]� ��������������������U��Q�M��M��E���E��t�M�Q��d�����E���]� ��������������������U��Q�M��EP�M�Q�rC������]� �������������������U��Q�M��E�P�~V������]����������U����M��E���	P�M��	Q�E@������~	�E�   ��E�    �E���]� ��������������������U��Q�M��EP�M�Q��������]� �������������������U��Q�M��E�����]����������������U���I���} t�^]����]����������U��Q����E��M����E���]���������������������U��   k� ǁ0��S�   �� ǂ0��N�   ��ǀ0�2k�   k�ǂ0�C_�   ��ǀ0��[�   k�ǂ0��S�   k�ǁ0��C�   k�ǀ0��j�   ��ǁ0��L�   k�	ǀ0�w:]���������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �}��   �/����u3���  ������u���3���  �j#���@�H���.������M����}��F���c��3��  ��/����|��,����|j �Z,������t��B���F���-��3��g  j� )�������������F  �} ��   �=�� ~{���������E�    �=� u�8���0��j��T8������ tj ������WK���GB���F������E������   ��} u�=|��t��E����3��   �   �}��   �|�R�{+�����E�}� uxh�   h �jh�  j��*�����E�}� tP�E�P�|�Q�;������t%j �U�R�(�����D�M��U��B�����j�E�P� ����3���3����}u
j �>a�����   �M�d�    Y_^[��]� ������������������������������������������������������������������������������������������������������������������������������������������������������������U��}u�>6���EP�MQ�UR�   ��]� ����������U��j�h8�h�Ld�    P���SVW���1E�3�P�E�d�    �e��E�   �} u�=�� u3��Z  �E�    �}t�}uT�=�� t�EP�MQ�UR����E�}� t�EP�MQ�UR�)���E�}� u�E�    �E������E���   �EP�MQ�UR�2���E�}u=�}� u7�EPj �MQ�z2���URj �EP�(���=�� t�MQj �UR����} t�}u@�EP�MQ�UR�(����u�E�    �}� t�=�� t�EP�MQ�UR����E��E������D�E���U܋E�P�M�Q�UR�EP�MQ�^����Ëe��E�    �E������E��
�E������E�M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������U��}u�EPj �MQ�h'���UR�EP������]�����������������������U��Qj j j���P�MQ�sI�����E��E���]�����������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_������������������������������������������������������������������������̀�@s�� s����Ë���������������������������̹   �-x���   �-����   �-x�f~�%���=  ��L  �Z���u���f/�v
�   �=  f/��!  �5p�f/��  fo�fs�fs���t:���f/�w,fW�f/�t"P��<$f�$f� Xu�   ��   3��   ��fW�f/���   �P��%X�fn-��fo���� fo�f��f��fs�4fo�f��fo�f��fo�f��fo�f��ff�fb�f��f��f��f��f��f��f��f��f~��� ~#f��f��f~�fs�f~��t
�   �    f~�fs�f~�ú   �   3��   �Ã� ��<$�$��t����u(�-���$�D$    �D$�D$�D$�9
���؃� ù   �-x���   �-����   �-x�fo�fs�f~�%���=  ��b���������fo�fs�fs����f/�v/��t�   �@����   �6�����   �*����   � ������f/�s'fW�f/��0����   ������   ���������fo؃�u�x�f/�rf\�fo�fs�#fs�#f~��t
�   ����f/�������p�f/������������u�*�����@��X��fn%��fn-��fn5��fn�fn�fb��    ��+�fn�f��fo�fs�3fs�3fo�fs�fs�ff�fb�f��ff�fb�f��f��fs�4f��Ë���;�u�*�Å��Y����=`��ك� ���E���V�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U������]�h��  h?  ��7�����E��E%�  =�  ��   ���E�$�2�����E��}�t�}�t!�}�t3�Jh��  �M�Q�7�����E�   h��  �U�R�7�����E���i�E�P���E�$j��0�����P�M�Q�E��s���$���E�$jj������&�U������U�E�E�h��  �M�Q�7�����E���]����������������������������������������������������������������������̃��$�B���   ��ÍT$���R��<$�D$tQf�<$t�I���   �u���=�� �O���   �����D���  �u,��� u%�|$ u���7���"��� u�|$ u�%   �t����-���   �=�� �����   ����(��Z�������������������������������������������������������U��E�<Ű� u�MQ�P������u
j������U�հ�P� ]��������������������U���!
����u�EPj �Hh�   �_/����]����������U����E�    �	�E����E��}�$}O�M��<Ͱ� t@�U��<մ�t3�E��Ű��M��U�R�j�E�P�������M��Ͱ�    ��E�    �	�U����U��}�$}3�E��<Ű� t$�M��<ʹ�u�U��հ��E�M�Q�뾋�]�����������������������������������������������������U��j�hX�h�Ld�    P���SVW���1E�3�P�E�d�    �E�   �=�� u�=D��j�..����h�   �.�����E�<Ű� t
�   �   h  h��jj� �����E�}� u�bJ���    3��jj
�������E�    �M�<Ͱ� u"j h�  �U�R�B2�����E�M�Ű��j�U�R�J�����E������   �j
��<����ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������U����E�    �E�    �	�E����E��}�$}F�M��<ʹ�u7kU������E��Ű��M����M�j h�  �U��հ�P�;1����뫸   ��]���������������������������������������������U��E�Ű�Q�]�����������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �e�} t8�E�8csm�u-�M�yu$�U�z �t�E�x!�t�M�y"�t�   �U�z ��   �E�H�y tS�E�    �U�B�HQ�U�BP�'���E������+�M��t	�E�   ��E�    �E�Ëe��]���E������,�U�B���t�U�B��M�}� t�U��M�Q�P�ҋM�d�    Y_^[��]���������������������������������������������������������������������������������U��Q�M��EP�M��?D���M����E���]� �����������U��Q�M��EP�M������M����E���]� �����������U��Q�M��E�� ��M�������]���������������������U��Q�M��M��<���E��t�M�Q�N�����E���]� ��������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �e�E�E��E�    �   k���E��M̋U�BP�M�Q������E���1�����   �U���1�����   �E���1���M���   ��1���U���   �E�    �E�   �E�   �E P�MQ�UR�EP�MQ�:@�����E��E�    ��   �U�R�  ��Ëe��m1��ǀ�      �E�H�MЋU�z�   �E�H���   �щU��	�E�H�MԋUԉU��E�H�M��E�    �	�U���U�E�M�;HsAkU��E؋M�;L~/kU��E؋M�;LkU��E؋L���M��U��EЋЉM��뫋U�R�EPj �MQ� �����E�    �E�    �E������E�    �   �   �   k���M�Ủ�E�P�{
�����f0���Mĉ��   �X0���U����   �E�8csm�u\�M�yuS�U�z �t�E�x!�t�M�y"�u/�}� u)�}� t#�U�BP�$3������t�M�Q�UR�5����ËE܋M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    PQSVW���3�P�E�d�    �e���.�����    u��.H���E�    � ����.���M���   j j �/���0)��E�������E������:����M�d�    Y_^[��]���������������������������������������������������U����E�E��}  t�M Q�UR�E�P�MQ��B�����}, u�UR�EP��;����MQ�U,R��;���E$�Q�UR�EP�M�Q��������U$�B���M�Ah   �U(R�E�HQ�UR�EP�M�Q�UR�f������E��}� t�EP�M�Q�)�����]����������������������������������������������������������U��Q�E��M��U��:csm�uN�E��xuE�M��y �t�U��z!�t�E��x"�u!�M��y u�-��ǀ�     �   ��3���]��������������������������������������U���D�E� �E� �E�x�   �M�Q���   �E��	�M�Q�U܋E܉E�}��|�M�U�;Q}���E���E�8csm��[  �M�y�N  �U�z �t�E�x!�t�M�y"��&  �U�z �  �6,�����    u�  �#,�����   �E�,�����   �M�E�j�UR�!������t��:E���E�8csm�u;�M�yu2�U�z �t�E�x!�t�M�y"�u�U�z u��D���+�����    ty�+�����   �E��+��ǀ�       �M�Q�UR�  ������t�C�M�Q�K  ���Ѕ�t+j�EP�����h$��M����h���M�Q��+��������U�:csm���  �E�x��  �M�y �t�U�z!�t�E�x"��i  �M�y �5  �U�R�E�P�M�Q�U R�EP�4�����E���M���M�U����U��E�;E���   �M��;U��E��M�;H~�˺   k� �M�A�E��U��B�E���M���M�U����U��}� ��   �E�H�Q���U��E�H�Q��E���M���M�U����U��}� ~d�E���MԋU�BP�M�Q�U�R��������u���E��E�P�M$Q�U R�E�P�M�Q�U�R�EP�MQ�UR�EP�MQ�P�����,�	���D���������(�U�%���=!�r���B���M�y t��B���U��tj�EP������M�����   �U�%���=!���   �M�y ��   �U�BP�MQ�/  ���Ѕ���   �)�����   �E���(�����   �M���(���U���   ��(���M���   �}$ u�UR�EP�6����MQ�U$R�6��j��EP�MQ�UR�������E�HQ�u������(���U���   �(���M���   �@�U�z v7�E��u*�M$Q�U R�E�P�MQ�UR�EP�MQ�UR�^  �� �������0(�����    u��kA����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���V�E�8  �u�o  ��&�����    tZ�&����j �9��   tC�M�9MOC�t8�U�:RCC�t-�E$P�M Q�UR�EP�MQ�UR�EP�&�������t�  �M�y t��?���U�R�E�P�MQ�U R�EP�0�����E���M����M��U����U��E�;E���   �M��U;|e�E��M;HZ�U��B�����M��Q�| t'�E��H�����U��B�L�   k� �L��u�U��B�����M��Q���@t�n���j�M$Q�U R�E�Pj �M��Q�����E�PR�MQ�UR�EP�MQ�UR������,�*���^��]������������������������������������������������������������������������������������������������������U����} t��)>���} u�h����E� �E�    �	�E����E��M�U�;}m�E�H�Q���U��E�H�Q��E���M���M�U����U��}� ~4�E���M�U�BP�M�Q�U����EPR�`������t�E���뀊E���]�����������������������������������������������U��Q�E�    �	�E����E��M�U�;}'h���E����M�Q�L�������t����2���]��������������������U��Q�#�����    t	�E�   ��E�    �E���]������������������������U����} t��<���E��M��}� t��<���U��:csm�u/�E��xu&�M��y �t�U��z!�t�E��x"�u��U<���M��Q�B���E�M��Q�B��M���U����U��E���E�}� ~0�M��U��E��H��Q�M���P��������u�   ��3���]�������������������������������������������������������������U��E�p�]����U��Q�E�M�M��U�z |'�E�H�U�
�M�Q�M��M��U�E�B�E��E���]���������������������������U��j�hؖh�Ld�    P���SVW���1E�3�P�E�d�    �e�E���   �t�U�U���E�H�U�D
�E��E�    �MQ�UR�EP�MQ�/�����E��}�t�}�t+�R�U��R�E�HQ������P�U�BP�M�Q������)j�U��R�E�HQ�����P�U�BP�M�Q��:���E�������   Ëe������E������M�d�    Y_^[��]�����������������������������������������������������������������������U��j�hx�h�Ld�    P���SVW���1E�3�P�E�d�    �e��E�    �E�x t-�M�Q�   k� �T
��t�E�x u�M���   �u3��j  �E���   �t�U�U���E�H�U�D
�E��E�    �M���   tn�E���td�=p� t[�p��E�j�U�R��������t6j�E�P��������t$�M�U܉�E��P�M�R������M����8���  �U���tXj�M�QR�������t9j�E�P�e������t'�M�U�B��M��Q�U�P������M���q8���@  �U���txj�M�QR�������tYj�E�P�������tG�M�QR�E�HQ�U�R�5������E�xu"�M�9 t�U��R�E�Q�;�����U����7���   �E�x uZj�M�QR�������t>j�E�P�������t,�M�QR�E��P�M�QR������P�E�P��������7���[j�M�QR�C������tAj�E�P�(������t/�M�QR�*������t�E���t	�E�   ��E�   ��,7���E�������   Ëe��_����E������E��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} u3��l�E��M��U��:csm�uW�E��xuN�M��y �t�U��z!�t�E��x"�u*�M��y u!����   �E��U�����M���   �3���]���������������������������������U���(�} u3���  �E��M��} t�   k� �M�T����   �E��8MOC�t�M��9RCC�t�U��@uz�E��8csm�uK�M��yuB�U��z �t�E��x!�t�M��y"�u�U��z u������    u3��H  ����   �E��E�����U��
�   �$  �E��8csm��  �M��y�  �U��z �t�E��x!�t�M��y"���   �U��z u#�.�����    u3���   ������   �E��M�M܋U�U؋E�   ��E؋M��Q�B���E�M��Q�B��M���U����U��E���E�}� ~d�M��U�E��HQ�U�R�E�P��������t?����   �E�M����E��} t�M�Q�U�R�EP�M�Q�
/�����   ��3���]����������������������������������������������������������������������������������������������������������������������������������������U��   ]�������U����E�    �E�E��   �� M��M��   �� U�U��} ��   �E�8 ��   �M��U��E��8csm�uD�M��yu;�U��z �t�E��x!�t�M��y"�u�U��z u�.�����   �E��M��QR�E�P�������E��
���M􋐈   ������M����   ������M����   ��U�������E�� ���������   �E�M����E�������    }���ǀ�       �   ��]���������������������������������������������������������������������������������������������U����E�E��   �� M��M��   �� U��U��E��8��G  �M�Q�������} ��   �������   �:csm�u~�������   �xum������   �y �t(������   �z!�t������   �x"�u1������   �QR�������tj�e�����   P�������Q�����   �9csm�um�>�����   �zu\�-�����   �x �t(������   �y!�t������   �z"�u �} t�����   �E�E����U�
�����M�����   �����M�����   ��]��������������������������������������������������������������������������������������������������U����E��M�U��E��}�RCC�t(�}�MOC�t�}�csm�t�@���ǀ�       ����������    ~�����   �E��M�����E��3��3���]����������������������������������������U��j�hx�h�Ld�    P���SVW���1E�3�P�E�d�    �e�E�x�   �M�Q���   �E��	�M�Q�U��E��E��J���   �E܋M܋���E܉�E�    �M�;M��   �}��~�U�E�;B}��U.���M�Q�E�M��E�   �U�B�M�|� t%�U�E؉Bh  �MQ�U�B�M�T�R�1���E�    ��E�P�!����Ëe��E�    �M؉M��f����E������   �)������    ~�s���   �EԋUԋ���MԉËU�;Uu��-���E�M�H�M�d�    Y_^[��]���������������������������������������������������������������������������������������������������U����E�     ������   �M��}� ��   �U��B�E��}� t%�M����t�E��H��U�E���E�M��R�U��B���E�M��Q��E���M����M��U���U�}� ~�E��M�U���t�M�   ���3���]������������������������������������������������U����������   u<�E�8csm�t1�M�9&  �t&�U�%���="�r�M�Q ��t
�   �  �E�H��ft4�U�z t�} uj��EP�MQ�UR�Y������   ��   ��   �E�x u$�M��������!���   �E�x ��   �M�9csm�uo�U�zrf�E�x"�vZ�M�Q�B�E��}� tH�M�Q�������t1�U$R�E P�MQ�UR�EP�MQ�UR�EP�U��� �E��E��7��+���)�M Q�UR�E$P�MQ�UR�EP�MQ�UR������ �   ��]���������������������������������������������������������������������������������������������������������U��Q�E�x t�M�Q�   k� �T
��u
�   �   �E���   t�U���t
�   �   �M�U�A;Bt$�M�Q��R�E�H��Q��������t3��O�U���t
�M���t1�E���t
�U���t�M���t
�E���t	�E�   ��E�    �E���]�������������������������������������������������������������U�������E��E��Hl�M��U�;4�t�E��Hp# �u����E��U����   ��]����������������������������U���]�������U��Q�}�   s	�E�   ��E�    �E���]�������������U��Q�EP�W*������u�M��_t	�E�    ��E�   �E���]����������������������������U��Q�EP�)������u�}_t	�E�    ��E�   �E���]����������������U��E��]������U����EP�M��L����M��)����t/�M��)����yt~�M��)��Ph  �UR�i������E��h  �EP�M��X)��P�������E��M��M��M��5����E���]����������������������������������U����EP�M������M���(����t/�M���(����yt~�M���(��Ph  �UR��������E��h  �EP�M��(��P�c������E��M��M��M������E���]����������������������������������U����EP�M������}	u	�E�@   �X�M��M(����t,�M��A(����yt~�M��1(��Pj@�UR�������E��j@�EP�M��(��P�������E��M��M��U��U�M�������E��]���������������������������������������������������U����EP�M��L����M��'����t,�M��'����yt~�M��'��Pj �UR�l������E��j �EP�M��^'��P�	������E��M��M��M��;����E���]����������������������������������������U��Q�EP�MQ���������u�}_t	�E�    ��E�   �E���]����������������������������U��Q�EP�MQ�:�������u�}_t	�E�    ��E�   �E���]����������������������������U����EP�M������M��\&����t,�M��P&����yt~�M��@&��Pj�UR�,������E��j�EP�M��&��P��������E��M��M��M�������E���]����������������������������������������U����EP�M��l����M��%����t/�M��%����yt~�M��%��Ph  �UR�������E��h  �EP�M��x%��P�#������E��M��M��M��U����E���]����������������������������������U����EP�M�������M��%����t,�M��%����yt~�M�� %��Pj�UR��������E��j�EP�M���$��P�������E��M��M��M������E���]����������������������������������������U����EP�M��,����M��|$����t/�M��p$����yt~�M��`$��PhW  �UR�I������E��hW  �EP�M��8$��P��������E��M��M��M������E���]����������������������������������U����EP�M������M���#����t,�M���#����yt~�M���#��Pj�UR�������E��j�EP�M��#��P�I������E��M��M��M��{����E���]����������������������������������������U����EP�M�������M��<#����t,�M��0#����yt~�M�� #��Pj�UR�������E��j�EP�M���"��P�������E��M��M��M�������E���]����������������������������������������U����EP�M��L����M��"����t,�M��"����yt~�M��"��Pj�UR�l������E��j�EP�M��^"��P�	������E��M��M��M��;����E���]����������������������������������������U����EP�M������M���!����t/�M���!����yt~�M���!��Ph�   �UR��������E��h�   �EP�M��!��P�c������E��M��M��M������E���]����������������������������������U��=4� uh  �EP�������j �MQ�=�����]����������������U��=4� uh  �EP�i������j �MQ������]����������������U��Q�=4� u'�}	u	�E�@   �j@�EP������E��E���j �MQ��������]���������������������������U��=4� uj �EP��������j �MQ�������]�������������������U��=4� uj�EP�������j �MQ�0�����]�������������������U��=4� uh  �EP�I������j �MQ�<�����]����������������U��=4� uj�EP�������j �MQ������]�������������������U��=4� uhW  �EP��������j �MQ�������]����������������U��=4� uj�EP�������j �MQ�������]�������������������U��=4� uj�EP�L������j �MQ������]�������������������U��=4� uj�EP�������j �MQ�"�����]�������������������U��=4� uh�   �EP��������j �MQ�B�����]����������������U��j j j�EP������]����������U����E�    �} u3��l�EP���������E��MQ�UR�EPj�M�Q�N������E��}� t5j jRh��hD�h`��UR�E�P�M�Q������P�s������E��3���]������������������������������������������U�������E��E��Hl�M��U�;4�t�E��Hp# �u�"���E��U��B��]�������������������������������U����6���E��E��Hl�M��U�;4�t�E��Hp# �u��
���E��U��B��]�������������������������������U��������E��E��Hl�M��U�;4�t�E��Hp# �u�b
���E��E��   ��]�����������������������������U����v���E��E��Hl�M��U�;4�t�E��Hp# �u�
���E��U��Bt��]�������������������������������U��Q�} u
����E���E��Qt�U��E���]�����������U���@���3ŉE��E�    �E�    �E�    �E�    �E�    �E�E��E�    �   ��U��
�    �-  �E�x u5�M��Qh  �   ��E���   Qj �U�R��������t�  j^h��jj�������E�jbh��jjh�  �m������E�jdh��jjh�  �R������E�jfh��jjh�  �7������E�jhh��jjh  �������Eԃ}� t�}� t�}� t�}� t�}� u��  �E��     �MԉM��E�    �	�U����U��}�   }�E�M���U���U��ۍE�P�M�QR�L��u�  �}�v�  �E�E�j �M�QRh�   �E��   Ph�   �Mԃ�Qh   �   ��E���   Qj �����$��u�?  j �U�BPh�   �M؁��   Qh�   �Uԃ�Rh   �   ���M���   Rj �l����$��u��  �}�~u�E�E��	�M���M�   k� �M����tQ�   �� �M����t>�   k� �U��
�E��	�M����M�   �� �E��9M��U�U�� ���j �E�HQ�U܁�   Rh   �E�Pjj �������u�E  �   k�3��M�f��   k��M�� �   k��M�� �   ���E�� �   ���U��
 �}�~�E�E��	�M���M�   k� �M����t[�   �� �M����tH�   k� �U��
�E��	�M����M�   �� �E��9M�� �  �E��M�f��A   ���h�   �U܁�   R�E�P�'�����j�MЁ�   Q�U�R������j�E�   P�M�Q��������U���    ��   �E���   �����J��   3�u#j hpjj h�   h��j�d�������u�j�U���   -�   P�������j�M���   ��   R�������j�E���   ��   Q������j�U���   P�������M��   �U�Ẻ��   �M܁�   �U���   �E��   �M���   �UЁ   �E���   �M؁��   �U���   �E�MȉHtj�U�R�0�����3���   j�E�P������j�M�Q������j�U�R�������j�E�P�������j�M�Q��������   �   �   �U���    tE�E���   �����Ju2�E���    w&hD�hpjj h�   h��j���������u̋Uǂ�       �Eǀ�       �Mǁ�   8��Uǂ�   ���Eǀ�   @��M�At   3��M�3��P�����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���,�} ~,�EP�MQ�  ���E�U�;U}�E���E��M�M�E�    �E�    �E�    �}$ u�U��H�M$�}( t	�E�	   ��E�   j j �UR�EP�M�Q�U$R��E��}� u3��<  �}� ~W3�uS�����3��u���rD�M���Q��������t#h��  �U��DP�O�����P�������E���E�    �M��M���E�    �U܉U�}� u3���  �E�P�M�Q�UR�EPj�M$Q���u
�  �z  j j �U�R�E�P�MQ�UR�p������E��}� u
�P  �K  �E%   tK�}  t@�M�;M ~
�.  �)  �U R�EP�M�Q�U�R�EP�MQ��������u
�   ��   ��   �U��U�}� ~W3�uS�����3��u��rD�M���Q�o�������t#h��  �U�DP�$�����P�������E���E�    �M؉M���E�    �UԉU��}� u�~�|�E�P�M�Q�U�R�E�P�MQ�UR�n�������u�V�T�}  u+j j j j �E�P�M�Qj �U$R��E��}� u�'�%�#j j �E P�MQ�U�R�E�Pj �M$Q��E��}� t�U�R��������E�P��������E���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�E��M�M��U��U�E����E��}� t�M����t�E����E��֋E+E�����]������������������������U��Q�E��;Ev	�E�   ��E�    �E���]�����������U��} t�E�M��U���U�E]������������������U����EP�M��L����M(Q�U$R�E P�MQ�UR�EP�MQ�UR�M��|��P�`�����$�E��M��_����E���]����������������������������U��Q�} t[�E���E�M��U��}���  u�EP�+�����3�}���  t*3�u&h��hpjj h  h��j���������u̋�]����������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�    �E�    �} ��   j j%hH�h��h��j"jh����EPj j �M�Q�Y�����P�f����� j&hL�jj�U�R�k������E܃}� u3���  j j)hH�h��h��j"jj��EP�M�Q�U�Rj �������P������ ��tj�E�P�9�����3��r  �M�Q�UR�b������E�j�E�P�������}� u3��D  �����E̋M̋Ql�UċE̋Hh�M��E�    j jEhH�h��h �j"j�U�Rj �E�Pj j �M�Q�O�����P�e����� ��t3���  jHhL�j�U���R�������E؃}� u3��  �   �� E؉E�j jOhH�h��h��j"j�M�Qj��U�R�E�P�M�Qj �������P������ ��tj�U�R������3��S  �EĉE�j�W������E�    �M���U�|
 t�E���M�| uC�U���E�| u�M���U�|
 t#hx�hpjj jYhH�j���������u̋M���U�|
 t/�E���M�T�����Huj�M���U�D
P�Z������M̋Qp��uI� ���u?�M���U�|
 t/�E���M�T�����Huj�M���U�D
P�������M؋U���M���U�E؉D
�M���U�EԉD
�E������   �j�q�����ËEԋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h �h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�   ��E�    �E��E܃}� u#hp�hpjj j6h��j覼������u̃}� u-�����    j j6h��h��hp��I�����3��  �} t	�E�   ��E�    �U؉Uԃ}� u#h�hpjj j7h��j�.�������u̃}� u-����    j j7h��h��h��������3��  �M���t	�E�   ��E�    �EЉẼ}� u#h0�hpjj j8h��j費������u̃}� u-����    j j8h��h��h0��U�����3��   �����E�}� u�����    3��t�E�    �U���u*����    �E�    j��M�Qh���_	�����E��9�U�R�EP�MQ�UR�w������E��E������   ��E�P�"�����ËEȋM�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������U��j@�EP�MQ������]����������U����} t	�E�   ��E�    �E��E��}� u&h`�hpjj h�   h��j�۹������u̃}� u0�0 ���    j h�   h��h��h`��{������   �-h�   �UR�EP��������M��U�: t3�������� ��]������������������������������������������������������������U����E�E��M��Q��   u�z����    ����   �E��H���U��J�}u�E�P�u ����E�E�E    �M�Q�V������U��B%�   t�M��Q����E��P�-�M��Q��t"�E��H��t�U��B%   u
�M��A   �UR�EP�M�Q�������P�W��������u	�E�������E�    �E���]����������������������������������������������������������������������U��j�h �h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h�hpjj jch��j荷������u̃}� u.������    j jch��h �h��0����������   �} t�}t�}t	�E�    ��E�   �U܉U؃}� u#h��hpjj jdh��j��������u̃}� u+�]����    j jdh��h �h������������H�MQ�������E�    �UR�EP�MQ�s������E��E������   ��UR�������ËEԋM�d�    Y_^[��]�����������������������������������������������������������������������������������������������������U��j@�EP�MQ������]����������U����} t	�E�   ��E�    �E��E��}� u&h`�hpjj h�   h��j諵������u̃}� u0� ����    j h�   h��h(�h`��K������   �-h�   �UR�EP�h������M��U�: t3������� ��]������������������������������������������������������������U��j�h@�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�   ��E�    �E��E܃}� u#hp�hpjj j6h��j膴������u̃}� u-������    j j6h��h�hp��)�����3��  �} t	�E�   ��E�    �U؉Uԃ}� u#h�hpjj j7h��j��������u̃}� u-�c����    j j7h��h�h�������3��  �M���t	�E�   ��E�    �EЉẼ}� u#h0�hpjj j8h��j蒳������u̃}� u-������    j j8h��h�h0��5�����3��   �i����E�}� u�����    3��t�E�    �U���u*�����    �E�    j��M�Qh���?�����E��9�U�R�EP�MQ�UR�������E��E������   ��E�P������ËEȋM�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������U����E�T=  �E�    �   k�����3���U�tj �E�P�U��E��}�zu�   �3���]���������������������U��Q�   k�����3���U�t�EP�U���]�������������������������U��Q�   k�����3���U�t�EP�U���]�������������������������U��Q�   k�����3���U�t�EP�MQ�UR�EP�U���MQ�U��R�E��P�MQ�`��]�������������������������������U��Q�   k�����3���U�t�EP�MQ�UR�EP�MQ�UR�U���EP�MQ�UR�EP����]�����������������������������U��Q�   k�����3���U�t�EP�MQ�UR�U��
jx�X2���]���������������������U��Q�   ������3���M�t�UR�EP�MQ�U��3���]�����������������������������U��Q�   k�����3���U�t�EP�MQ�UR�U��3���]�����������������������������U��Q�   k� ����3���U�t	�EP�U���p��]�����������������U��Q�   �� ����3���M�t	�UR�U��
�EP�|��]�����������������������������U��Q�   ������3���M�t	�UR�U��
�EP�t��]��������������U��Q�   k�����3���U�t�EP�MQ�U���UR�EP�x��]���������������������U��Q�   k�����3���U�t�U���]�������������U��Q�   ������3���M�t�UR�EP�U���]���������������������U��Q�   k�����3���U�t�U��3���]�������������������������U��Q�   k�����3���U�t�EP�MQ�UR�EP�U��
jx�X3���]�����������������U��Q�   k�����3���U�t�EP�MQ�U��
jx�X3���]�������������������������U���H�E�P���M��t	�U�U���E�
   f�E���]�����������������U��Q�   k�����3���U�t�U����3ҋ�]�������������������U��Q�   ������3���M�t�UR�EP�MQ�U���UR�EP�\�   ��]����������������������������U��Q�=� }
��������=� ~	�E�   ��E�    �E���]��������������������������U��Qh@����E�h`��E�P��3���   k� ����hl��E�P��3���   �� ����hx��U�R��3���   �ቁ��h���U�R��3���   k�����h���E�P��3���   ������h���U�R��3���   k�����h���E�P��3���   k�����h���E�P��3���   k�����h��E�P��3���   ������h ��U�R��3���   k�	����h8��E�P��3���   k�
����h`��E�P��3���   k�����h|��E�P��3���   k�����h���E�P��3���   k�����h���E�P��3���   k�����h���E�P��3���   k�����h���E�P��3���   ������h��U�R��3���   k�����h0��E�P��3���   k�����hX��E�P��3���   k�����hp��E�P��3���   k�����h���E�P��3���   k�����h���E�P��3���   k�����h���E�P��3���   k�����h���E�P��3���   k�����h���E�P��3���   k�����h���E�P��3���   k�����h��E�P��3���   k�����h0��E�P��3���   k�����h@��E�P��3���   k�����hX��E�P��3���   k�����hl��E�P��3���   k�����h���E�P��3���   ��������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�   ������3���M�t�UR�EP�MQ�UR�U��
jx�X3���]�����������������U��Q�   k�����3���U�t	�EP�U��3���]���������������������U��Q�   k�	����3���U�t�EP�MQ�UR�EP�U���]�����������������������������U��Q�   k�����3���U�t�EP�MQ�UR�U���]�����������������U��EP�T]������������������U��EP�d]������������������U��EP�hP�l]�����������U��j �T�EP�P]����������U��Q�   k�
����3���U�t�EP�MQ�U���]���������������������U��Q���E��M��#M��U#Uʉ��E���]������������������������U��Q�E�    ����t
j
�����������E��}� t
j�Ǳ��������t#j�������t�   �)jh  @j�V�����j葥����]���������������������������������U���Ph��  h?  �*������E��E%�  =�  ��   ���E�$��������E��}� ~R�}�~�}�t�Dh��  �M�Q��������E�j  �U�R�E�]��E؃��$���E�$j�+������?  �E�P�E��s���$�E�]��EЃ��$���E�$jj�ɡ����$�  �E��������Dzh��  �M�Q�L������E��  �U�R���E�$�������]�} }!�   �+E9E�}	�E�   ��	�M�M�M������+U9U�~	�E�����	�E�E�E��}� 
  ~M�M�Q���E��$���p��$�`������$�E�]��Eȃ��$���E�$jj������$�(  �}�   ~T�U���   R���E��$�������]��E�P���E��$�E�]��E����$���E�$jj葠����$��   �}����}<�M�Q�E���s���$�E�]��E����$���E�$jj�L�����$�   �}����}Q�U���   R���E��$�c������]��E�P���E��$�E�]��E����$���E�$jj������$�,�M�Q���E��$�������]�h��  �U�R�k������E���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�E��M�Q�UR�ӱ������]�������������������U��Q�E�E��M�Q�UR�EP��������]���������������U��Q�E�E��M�Q�UR��������]�������������������U��Q�E�E��M�Q�UR�EP��������]���������������U��Q�E�E��M�Qj �UR�EP�MQ�UR�.�������]���������������������U��Q�E�E��M�Q�UR�EP�MQ�UR�EP���������]�������������������U��Q�E�E��M�Q�UR�EP�MQ���������]�����������U��Q�E�E��M�Qj �UR�EP�MQ�G�������]�������������������������U��Q�E�E��M�Q�UR�EP�MQ�UR��������]�����������������������U��Q�E�E��M�Q�UR�EP�MQ�UR��������]�����������������������U���D�E�    3��E��EĉEȉẺEЉEԉE؍M��M��} t	�E�   ��E�    �U��U�}� u#h��hpjj jih��j�*�������u̃}� u.�����    j jih��hD�h�������������  �} t	�E�   ��E�    �M��M�}� u#hX�hpjj jnh��j豜������u̃}� u.�����    j jnh��hD�hX��T���������   �E�E��M��A����U��BB   �E��M�H�U��E��M�Qj �UR�E�P�S������E�} u�E��Q�M��Q���U�E��M�H�}� |"�U���  3Ɂ��   �M܋U�����M����U�Rj �/������E܋E��]�����������������������������������������������������������������������������������������������������������������U��Q�E�E��M�Qj �UR�EP�MQ�C�������]������������������������̋T$�L$��   u@�:u2��t&:au)��t��:Au��t:au������uҋ�3���������Ë���   t���:u����t���   t�f���:u΄�t�:auń�t����������������������������������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^����������������������������U����F����E��E��Hl�M��U�;4�t�E��Hp# �u������E�� ���]��������������������������������U��Q�����E��}� u	������E�����]������������U��V�Ǟ���M��UR�d�������������0^]�����������U��Q�����E��}� u	������E�����]������������U����} t	�E�   ��E�    �E��E��}� u&h��hpjj h�   h��j�ۘ������u̃}� u%j h�   h��h �h���������   ������U� �3���]��������������������������������������U����} t	�E�   ��E�    �E��E��}� u&h��hpjj h�   h��j�+�������u̃}� u%j h�   h��h�h����������   ��[����U� �3���]��������������������������������������U��Q�E�    �	�E����E��}�-s�M��U;͐�u�E��Ŕ��7�ԃ}r�}$w	�   �"� �}�   r�}�   w	�   ���   ��]�������������������������������U��Q�����E��}� u	�   ���`����M�3���]����������������������U��Q�V����E��}� u	�   ���9����M�3���]����������������������U��j�hd�    P�����3�P�E�d�    �EP�M��M����E�    �M�M�M������P�E�L#Mu;�} t�M��q�������   �M�H#U�U���E�    �}� u	�E�    ��E�   �E�E��E������M������E�M�d�    Y��]�������������������������������������������������U��jh  �EPj �������]�������U��jh  �EP�MQ�������]���������������������U��jh  �EPj ������]�������U��jh  �EP�MQ������]���������������������U��Q�}	u	�E�@   �jj@�EPj �N������E��E���]������������������U��Q�}	u	�E�@   �jj@�EP�MQ�������E��E���]����������������U��jh  �EPj �������]�������U��jh  �EP�MQ������]���������������������U��jj �EPj ������]����������U��jj �EP�MQ�l�����]��������U��j �EP������]��������������U����EP�M�謝���M�������x t8�M�������H�y�  u$jj �UR�EP��������E��M�躭���E���E�    �M�覭���E���]�����������������������������������U��jj �EPj ������]����������U��jj �EP�MQ�|�����]��������U��jj �EPj �^�����]����������U��jj �EP�MQ�<�����]��������U��jj �EPj ������]����������U��jj �EP�MQ�������]��������U��jhW  �EPj �������]�������U��jhW  �EP�MQ������]���������������������U��jj�EPj ������]����������U��jj�EP�MQ�l�����]��������U��jj �EPj �N�����]����������U��jj �EP�MQ�,�����]��������U����E�E��M���U��E����E��}� t��E�+E������]����������������������������U��j �������]������������������U���(V�E�    �EP�M������M��d�������   �U��E�    �	�E����E��}�s3�M��U��P�2��������M��U�D�P������E�L0�M��jChD�j�U��R�������E��}� ��   �E��E��E�    �	�M����M��}���   �U��:�E����E�j jJhx�h��h���M��U��P�M���U�+U�+�Q�E�P�������P�0������M�Q�n�����E��E��U��:�E����E�j jMhx�h��hx��M��U�D�P�M���U�+U�+�Q�E�P������P�͚�����M�Q������E��E��#����U�� �E����E��M��M�M��ש���E�^��]�������������������������������������������������������������������������������������������������������������������U��j 褙����]������������������U���(V�E�    �EP�M��Ԙ���M��$�������   �U��E�    �	�E����E��}�s4�M��U�D�8P���������M��U�D�hP�ܸ����E�L0�M��jjhD�j�U��R蠊�����E��}� ��   �E��E��E�    �	�M����M��}���   �U��:�E����E�j jqhx�h��h��M��U�D�8P�M���U�+U�+�Q�E�P������P�������M�Q�,�����E��E��U��:�E����E�j jthx�h��h���M��U�D�hP�M���U�+U�+�Q�E�P�W�����P苘�����M�Q�ɷ����E��E��"����U�� �E����E��M��M�M�蕧���E�^��]�����������������������������������������������������������������������������������������������������������������U��j �������]������������������U��j �EP�MQ�UR�EP�MQ������]��������������U���T�E�    �E�    �E�    �EP�M��W����} t	�E�   ��E�    �M�M�}� u&h��hpjj h�   hx�j�J�������u̃}� u@�����    j h�   hx�h(�h����������E�    �M�� ����E��  �} t	�E�   ��E�    �E�E��}� u&hD�hpjj h�   hx�j輋������u̃}� u@�����    j h�   hx�h(�hD��\������E�    �M�蒥���E��  �U� �} t	�E�   ��E�    �E܉E؃}� u&hl�hpjj h�   hx�j�(�������u̃}� u@�}����    j h�   hx�h(�hl���������E�    �M�������E���  �} t	�E�   ��E�    �UԉUЃ}� u&h��hpjj h   hx�j蚊������u̃}� u@������    j h   hx�h(�h���:������E�    �M��p����E��^  j j j��MQj �M��]�����BP��E��}� u��P���������   h
  hD�j�M���Q�������E��}� u��   �U�R�E�Pj��MQj �M��������BP���u��P�|������   h  hD�j�M��Q衅�����E��}� u�k�UR�EP�MQ�U�R�EP�M�Q�������E�}� tBj j �UR�EPj��M�Qj �M��f�����BP���u��P�������E�    j�M�Q赗����j�U�R觗�����E�E��M������E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP�MQ�/�����]��������������U��j j �EP�MQ�UR�EP������]����������������U���   V�E�E��M����M��}�v��  �U������$�8��M�y |�U�zǅl���   �
ǅl���    ��l����E�}� u&h�hpjj h�  h �j��������u̃}� u0�\����    j h�  h �h,h�������3��X  �UR�EP�M�Q�E����   Q�  ���-  �U�z |�E�x	�E�   ��E�    �M��M܃}� u&h�hpjj h�  h �j�W�������u̃}� u0�����    j h�  h �h,h��������3��  �EP�MQ�U�B�M����   R�j  ���}  �E�x |�M�yǅ\���   �
ǅ\���    ��\����Uԃ}� u&hPhpjj h�  h �j螅������u̃}� u0������    j h�  h �h,hP�>�����3���  �MQ�UR�E�H�U����   P�  ����  �M�y |�U�z	�E�   ��E�    �E��Ẽ}� u&hPhpjj h�  h �j��������u̃}� u0�C����    j h�  h �h,hP������3��?  �UR�EP�M�Q�E���  Q�  ���  �}  ��   �UR�EP�MQ�URj�EP�4  ����u3���  �M�9 u3���  �U��    f��U����M��U����M��UR�EP�MQ�URj�EP��  ����u3��  �   �MQ�UR�EP�MQj �UR�  ����u3��Y  �E�8 u3��J  �M��    f��M����E��M����E��MQ�UR�EP�MQj�UR�H  ����u3���  ��  �E�x|�M�yǅt���   �
ǅt���    ��t����Uă}� u&h�hpjj h(  h �j��������u̃}� u0�f����    j h(  h �h,h�������3��b  �M Q�UR�EPj�M�QR�h  ���;  �E�x |�M�y	�E�   ��E�    �U��U��}� u&hhhpjj h1  h �j�e�������u̃}� u0�����    j h1  h �h,hh������3��
  �M Q�UR�EPj�M�QR�  ���
  �E�x |�M�yǅd���   �
ǅd���    ��d����U��}� u&hhhpjj h9  h �j谁������u̃}� u0�����    j h9  h �h,hh�P�����3��
  �M�A��   ���U��}� u�E�   �U R�EP�MQj�U�R��  ���	  �E�x |�M�ym  	�E�   ��E�    �U��U��}� u&h�hpjj hD  h �j��������u̃}� u0�;����    j hD  h �h,h�膿����3��7	  �M Q�UR�EPj�M�Q��R�:  ���	  �E�x |�M�y	�E�   ��E�    �U�U��}� u&hPhpjj hM  h �j�7�������u̃}� u0�����    j hM  h �h,hP�׾����3��  �M Q�UR�EPj�M�Q��R�  ���^  �E�x |�M�y;ǅ|���   �
ǅ|���    ��|����U�}� u&h�hpjj hV  h �j�������u̃}� u0������    j hV  h �h,h�������3���  �M Q�UR�EPj�M�QR��  ���  �E�x |�M�y	�E�   ��E�    �U��U؃}� u&hhhpjj h^  h �j��~������u̃}� u0�(����    j h^  h �h,hh�s�����3��$  �M�y%�UR�EP�   k� �E��L  Q��  ���#�UR�EP�   �� �U��
L  P�  ����  �M�9 |�U�:;	�E�   ��E�    �EЉEȃ}� u&hhpjj hi  h �j��}������u̃}� u0�J����    j hi  h �h,h蕼����3��F  �U R�EP�MQj�U�P�M  ���   �M�y |�U�z	�E�   ��E�    �E��E��}� u&h�hpjj hp  h �j�J}������u̃}� u0�����    j hp  h �h,h�������3��  �U�B�E��Y  �T  �M�y |�U�z	�E�   ��E�    �E��E��}� u&h�hpjj hw  h �j�|������u̃}� u0�����    j hw  h �h,h��M�����3���  �U R�EP�MQj�U�BP�
  ����  �M�y |�U�z	�E�   ��E�    �E��E��}� u&h�hpjj h~  h �j�|������u̃}� u0�V����    j h~  h �h,h�衺����3��R  �U�z u	�E�   ��E�H���M�U�z |�E�xm  	�E�   ��E�    �M��M��}� u&h�hpjj h�  h �j�V{������u̃}� u0�����    j h�  h �h,h��������3��  �E�H;M�}	�E�    �-�U�B��   ���E��U�B��   ��;U�|	�U����U��E P�MQ�URj�E�P�o  ���B  �}  t+�MQ�UR�EP�MQj�UR�f
  ����u3��  �)�EP�MQ�UR�EPj �MQ�;
  ����u3���  ��  �UR�EP�MQ�URj�EP�
  ����u3��  �  �M�y |	�E�   ��E�    �U���x�����x��� u&h�hpjj h�  h �j��y������u̃�x��� u0�4����    j h�  h �h,h�������3��0  �M�A��d   ���U��U R�EP�MQj�U�R�(  ����  �E�x����|�M�y�  ǅp���   �
ǅp���    ��p�����h�����h��� u&h�hpjj h�  h �j�y������u̃�h��� u0�b����    j h�  h �h,h�護����3��^  �M�A��d   ����k�d�U�B��d   ��ʉM��E P�MQ�URj�E�P�@  ���  �����E�    �M�y  tǅ`���   �
ǅ`���    j h�  h �h,hpj"j�URj�諠����`�����R�E�Q�U�P�M�Q������P�ru���� ��X�����X���Pu�U�    ��E����M�+ЋE��M��E��LB��U�
�Y�E��%   f��E����U�
�E����U�
�0�.3�u&hhhpjj h�  h �j�w������u�3���   ^��]ÍI ��ҭ��g����ͥb��T�H�0��E����;�l�������v���  	
���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �} t�EP�MQ�UR�   ���   �E�M;sn�U���U�	�E���E�M��t3�E��
   ����0�E��Ef�A�E��
   ���E�U����U�뼋E��U��Q�M��U�+E��M��	�U�    ��]��������������������������������������������������U����E��M��U�:vF�E��
   ����0�E�f��M����M��U����M��E��
   ���E�} ~�U�:w��E��M�U�E���M����M��U�f�f�E��M��U�f�f��M����M��U�f�E�f��M���M�U�;U�rƋ�]����������������������������������������������U��E�8 t=�M���t3�E��Uf�f��M����E��M���M�U����M��]�����������������������U���h���3ŉE��E�E��}� t�}�t��M��T  �U���E��X  �M���U��\  �E�M���   ��  �E�   �}t�E�    �U�Bl  f�E�M�Q��f�U�Ef�Hf�M�Uf�Bf�E�Mf�Qf�U��Ef�f�M�3�f�U��}� t%j j �E�P�M�Qj �U��`  P�������E��#j j �M�Q�U�Rj �E��`  Q�̯�����E؃}� �  �U���R�|{������t#h��  �E؍L Q�1�����P�԰�����E���E�    �U��Ũ}� ��   �}� t)�E�P�M�Q�U�R�E�Pj �M��`  R�^������E��'�E�P�M�Q�U�R�E�Pj �M��`  R� ������E؋ẺE܋M؃��M؃}� ~;�U�: v3�E��U�f�f��M����E��M܃��M܋U����M�붋U�R�������   �  �E������  �U�: ��  3�f�E��E�    �E�    �M�M��	�U����U��E���M��U���E��M܃��M܋U�;U�u�ҋE܃��E܋M���UċEă�'�Eă}�R�
  �M���Ի�$����E��E��M����M��}�w0�U��$�(��E�   �m   f�E���b   f�M��	�B   f�U��  �E��EȋMȃ��Mȃ}�w0�U��$�8��E�   �d   f�E���a   f�M��	�A   f�U��e  �E��E��}�t�}�t��y   f�M��	�Y   f�U��8  �E��E��}�t�}�t	��E�   �I   f�M��  �U��U��}�t�}�t	��E�   �H   f�E���  �M��M��}�t�}�t	��E�   �M   f�U��  �E��E��}�t�}�t	��E�   �S   f�M��  h��U�R�J�������u�E��
�E��h��M�Q�*�������u	�U���Uܸp   f�E��H  �M�y�   k� �M��L  �U���   �� �M��L  �Uԃ}�u;�E�8 v3�M��E�f�f�
�U����M��Uԃ��UԋE����U�
�E�E����t;�U�: v3�E��U�f�f��M����E��Mԃ��MԋU����M�뻋U܉U�������E���ti�M��U�J�E�M����tQ�E�8 tI�M����'u�E���E��3�M��E�f�f�
�U����M��U���U�E����U�
���E��M�A�U��m����E��t5�M�Q�UR�EP�MQ�UR�E�P�MQ���������u3��C�U܉U��1�E��U�f�f��M����E��M���M�U����M�������   �M�3��ˈ����]Ë������'�q��:�c�ع�� � 







































































	�F�M�X�c�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j ��~����]������������������U���(V�E�    �EP�M��4q���M�脴������   �U��E�    �	�E����E��}�s:�M��U싄��   P�֐�������M��U싄��   P辐����E�L0�M��jHh��j�U�DP��b�����E��}� �  �M��M��E�    �	�U����U��}���   �:   �M�f��U����U�j jOh �hd�h���E��M싔��   R�E���M�+M���+�P�U�R読����P�=q�����E�P�������M��A�U��:   �M�f��U����U�j jRh �hd�h �E��M싔��   R�E���M�+M���+�P�U�R�:�����P��p�����E�P蓏�����M��A�U�����3��M�f��U����U��E��E�M������E�^��]������������������������������������������������������������������������������������������������������������������������������U��j �#m����]������������������U���(V�E�    �EP�M���n���M���������   �U��E�    �	�E����E��}�s:�M��U싄��   P�f��������M��U싄�  P�N�����E�L0�M��joh��j�U�DP�`�����E��}� �  �M��M��E�    �	�U����U��}���   �:   �M�f��U����U�j jvh �h� h� �E��M싔��   R�E���M�+M���+�P�U�R�:�����P��n�����E�P蓍�����M��A�U��:   �M�f��U����U�j jyh �h� h8�E��M싔�  R�E���M�+M���+�P�U�R�ʪ����P�]n�����E�P�#������M��A�U�����3��M�f��U����U��E��E�M��b}���E�^��]������������������������������������������������������������������������������������������������������������������������������U��j �h����]������������������U���T�EP�M��\l���M�謯������   �U��E�    �E�d  �E�    �E�    �	�E����E��}���  �}�uWh�   h��j�M�Q�=^�����E��}� u�E�    �M��1|���E��  �U�Rj �E�P�������M��M��E�d  �E�    �	�U���U�}���   �E�3ҹ   ���t�U����U���}�uQ�E�E��M�U���j h�   h �h�h��E�M��R�E�+E�P�M�U���P�
�����P�>l�����M�U��P�v������M��T�U��Z����E�    �	�E���E�}���   �E�3ҹ   ���t�U����U���}�uT�E�E��M�U��D�j h�   h �h�h��E�M�T�R�E�+E�P�M�U��D�P�X�����P�k�����M�U�D�P�Ê�����M��T�U��V����E�    �	�E����E��}���   �E�3ҹ   ���t�U����U���}�uT�E�E��M��U��D�8j h�   h �h�hp�E��M�T�8R�E�+E�P�M��U��D�8P襧����P��j�����M��U�D�8P�������M��T�U��V����E�    �	�E܃��E܃}���   �E�3ҹ   ���t�U����U���}�uT�E�E��M܋U��D�hj h�   h �h�hP�E܋M�T�hR�E�+E�P�M܋U��D�hP������P�&j�����M܋U�D�hP�]������M��T�U��V����E�    �	�E؃��E؃}���   �E�3ҹ   ���t�U����U���}�u]�E�E��M؋U�����   j h�   h �h�h�E؋M􋔁�   R�E�+E�P�M؋U�����   P�6�����P�ji�����M؋U􋄊�   P螈�����M��T�U��J����E�3ҹ   ���t�U����U���}�uQ�E�E��M����   j h�   h �h�h��U􋂠   P�M�+M�Q�U����   P蟥����P��h�����M􋑠   R�������M��T�U��E�3ҹ   ���t�U����U���}�uQ�E�E��M����   j h�   h �h�h��U􋂤   P�M�+M�Q�U����   P������P�Eh�����M􋑤   R�}������M��T�U��E�3ҹ   ���t�U����U���}�uQ�E�E��M����   j h�   h �h�hx�U􋂨   P�M�+M�Q�U����   P胤����P�g�����M􋑨   R�������M��T�U��}�u�E��M􋑬   ���   �E�ǀ�       �E�    �	�Mԃ��Mԃ}���   �E�3ҹ   ���t�U����U���}�ud�E���M��A�EԋM�����   j h�   h �h�h@�UԋE􋌐�   Q�U�+U���R�EԋM�����   R�B�����P��f�����EԋM􋔁�   R葅�����M��TA�U��C����E�    �	�EЃ��EЃ}���   �E�3ҹ   ���t�U����U���}�ud�E���M��A�EЋM�����   j h�   h �h�h0	�UЋE􋌐�   Q�U�+U���R�EЋM�����   R�|�����P�f�����EЋM􋔁�   R�˄�����M��TA�U��C����E�    �	�Ẽ��Ẽ}���   �E�3ҹ   ���t�U����U���}�ud�E���M��A�E̋M�����   j h�   h �h�h
�ŰE􋌐�   Q�U�+U���R�E̋M�����   R趡����P�Ie�����E̋M􋔁�   R�������M��TA�U��C����E�    �	�Eȃ��Eȃ}���   �E�3ҹ   ���t�U����U���}�ud�E���M��A�EȋM����  j h�   h �h�h �UȋE􋌐  Q�U�+U���R�EȋM����  R������P�d�����EȋM􋔁  R�?������M��TA�U��C����E�    �	�Eă��Eă}���   �E�3ҹ   ���t�U����U���}�ud�E���M��A�EċM����L  j h�   h �h�h��UċE􋌐L  Q�U�+U���R�EċM����L  R�*�����P�c�����EċM􋔁L  R�y������M��TA�U��C����E�3ҹ   ���t�U����U���}�uX�E���M��A�E���T  j h�   h �h�h��M�T  R�E�+E���P�M���T  R茟����P�c�����E�T  Q�߁�����U��DB�E��E�3ҹ   ���t�U����U���}�uX�E���M��A�E���X  j h�   h �h�h��M�X  R�E�+E���P�M���X  R�������P�b�����E�X  Q�J������U��DB�E��E�3ҹ   ���t�U����U���}�uX�E���M��A�E���\  j h�   h �h�hx�M�\  R�E�+E���P�M���\  R�b�����P��a�����E�\  Q赀�����U��DB�E��E�3ҹ   ���t�U����U���}�uX�E���M��A�E���`  j h�   h �h�hX�M�`  R�E�+E���P�M���`  R�͝����P�`a�����E�`  Q� ������U��DB�E������M��M��M��op���E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�EP�MQ�n����]��������������U���l�E�    �E�E��MQ�M��\���} t	�E�   ��E�    �U�U��}� u&h��hpjj h  h �j�R������u̃}� u@������    j h  h �hHh���B������E�    �M��xl���E��  �} t	�E�   ��E�    �M�M�}� u&hD�hpjj h  h �j�R������u̃}� u@�i����    j h  h �hHhD�贐�����E�    �M���k���E��   3��Mf��} t	�E�   ��E�    �U�U��}� u&hl�hpjj h  h �j�~Q������u̃}� u@�ӗ���    j h  h �hHhl��������E�    �M��Tk���E��j  �} u�M��G�������   �U���E�E܋M܉M��U�U��}� �N  �E��M؃}� t�}�%t
�  �/  �} t	�E�   ��E�    �UԉUЃ}� u&hdhpjj h7  h �j�P������u̃}� u@�����    j h7  h �hHhd�:������E�    �M��pj���E��  �M���M�E�    �U���#u�E�   �M���M�U�R�E�P�M�Q�UR�EP�M�R�M��#���P�g�������u�}� v�E�   �7�E���E�'�M�Uf�f��M���M�U���U�E����E������}� u,�}� v&3ɋUf�
�E+E��E��M��i���E��   �   3ɋU�f�
�}� u�}� w�ȕ��� "   �v�E�    �}� u&h�hpjj hw  h �j�-O������u̃}� u=肕���    j hw  h �hHh��͍�����E�    �M��i���E���E�    �M���h���E���M���h����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP�MQ�i����]��������������U��j j �EP�MQ�UR�EP��h����]����������������U��E�� ]������U���<�EP�M���V���}   ��   �M��?�����t,�M��3�����yt~�M��#���Pj�UR�a�����E��j�EP�M�����P�H�����E��}� t,�M���������   �E��M�M���f���E��  ��U�U��M��f���E��  �M�襙��� �xt~q�M�蕙��P�M�����   Q蟚������tO�U�����   �   k� �T��   �� �E�D��   ��M�}�s������U��D� �E�   �=�j���� *   �   k� �U�T��E�   �}�s�貊���E��D� �E�   j�M�������QRj�E�P�M�Q�U�Rh   �M��Ę��� �   �ዔ�   R�M�諘��P�n�����$�E�}� u�E�E܍M��e���E��\�}�u�   k� �D��E؍M��_e���E��9�/�   �� �T��   k� �D���ЉUԍM��.e���E���M��!e����]�������������������������������������������������������������������������������������������������������������������������������������������������U��Q�=4� u$�}A|�}Z�E�� �E���M�M��E���j �UR�.s������]�����������������������������̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[����������������������������������������������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ����������������������������������������U����E�E��M�M��U���M��+�P�  ����]��������������������U��� �E�E��M�M�U�E��
;��   �U�U��E�E�M�Q�U�R�������E��}� t�E��E��s�M���Q�U��R�^������E��}� t�E��E��F�M���Q�U��R�7������E��}� t�E��E���M���Q�U��R�������E��E��E�M�M�E��3���]����������������������������������������������������U��Q�} t�} ~	�E�   ��E������E��E�E��]��������������������U����E�E�M�M�U���M��;�tK�E�E��M�M�U�R�E�P�E������E��}� t�M��M���U���R�E��P�������E��E��3���]������������������������������U���(�E�E��M�M�U�U��}��g  �E��$����M�Q�U�R�������E��}� t�E��E��s�M���Q�U��R�������E��}� t�E��E��F�M���Q�U��R�i������E��}� t�E��E���M���Q�U��R�B������E�E�E�M�M�E���   �U�R�E�P�������E��}� t�M��M��F�U���R�E��P��������E��}� t�M��M���U���R�E��P��������E��M��M܋E��i�U�R�E�P�������E��}� t�M��M���U���R�E��P�������E؋E��*�M�Q�U�R�p������3���EP�M�Q�U�R�   ����]ÍI ����D���<�������������������������������������������������������������������������������������������������������������������������U����} �R  �EP�MQ��������E��}� t�E��O  �U��R�E��P�������E��}� t�E��(  �M��Q�U��R�������E��}� t�E��  �E��P�M��Q�n������E��}� t�E���  �U��R�E��P�G������E��}� t�E��  �M��Q�U��R� ������E��}� t�E��  �E��P�M��Q��������E��}� t�E��e  �U��R�E��P��������E��}� t�E��>  �M�� �M�U�� �U�E�� �E�����MM�M�UU�U�E�E��}���  �M��$����U��R�E��P�_������E��}� t�E���  �M��Q�U��R�8������E��}� t�E��  �E��P�M��Q�������E��}� t�E��}  �U��R�E��P��������E��}� t�E��V  �M��Q�U��R��������E��}� t�E��/  �E��P�M��Q�������E��}� t�E��  �U��R�E��P�u������E��}� t�E���  3���  �M��Q�U��R�G������E��}� t�E��  �E��P�M��Q� ������E��}� t�E��  �U��R�E��P��������E��}� t�E��e  �M��Q�U��R��������E��}� t�E��>  �E��P�M��Q�������E��}� t�E��  �U��	R�E��	P�������E��}� t�E���  �M��Q�U��R�]������E��}� t�E���  �E��P�M��Q��������  �U��R�E��P�������E��}� t�E��  �M��Q�U��R��������E��}� t�E��`  �E��P�M��Q��������E��}� t�E��9  �U��R�E��P�������E��}� t�E��  �M��Q�U��R�������E��}� t�E���  �E��
P�M��
Q�X������E��}� t�E���  �U��R�E��P�1������E��}� t�E��  �M��Q�U��R�J������  �E��P�M��Q��������E��}� t�E��[  �U��R�E��P��������E��}� t�E��4  �M��Q�U��R�������E��}� t�E��  �E��P�M��Q�z������E��}� t�E���   �U��R�E��P�S������E��}� t�E��   �M��Q�U��R�,������E��}� t�E��   �E��P�M��Q�������E��}� t�E��t�U��R�E��P�������E��}� t�M��M��F�U��R�E��P�z������E��}� t�M��M���U��R�E��P�S������E�M�M��E��3���]�����#�L�������(��������j�������C�[������4�`������9�e������>�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���@���3ŉE��} ~�EP�MQ��  ���E��}�}3���  �}  ~�U R�EP��  ���E ��} �}3��  �E�    �}$ u�M��B�E$�} t
�}  ��  �M;M u
�   �o  �} ~
�   �_  �}~
�   �O  �U�R�E$P�L��u3��6  �} u�} t2�}u�}  t&h�hpjj h�   hpj�:������u̃} ��   �}�s
�   ��  �U�U��	�E���E�   k� �E����tQ�   �� �E����t>�U��   k� �M��;�|#�E��   �� �E��;�
�   �k  듸   �_  �}  ��   �}�s
�   �E  �E�E��	�M���M�   k� �M����tQ�   �� �M����t>�E��   k� �U��;�|#�M��   �� �M��;�
�   ��  듸   ��  j j �MQ�URj	�E$P��E��}� u3��  �}� ~W3�uS�����3��u���rD�U���R�mE������t#h��  �E��L Q�"c����P��z�����E���E�    �UЉU���E�    �E��E؃}� u3��'  �M�Q�U�R�EP�MQj�U$R���u
��   ��   j j �E P�MQj	�U$R��E܃}� u
��   ��   �}� ~W3�uS�����3��u܃�rD�M���Q�D������t#h��  �U܍DP�Vb����P��y�����E���E�    �MĉM���E�    �ỦUԃ}� u�Q�O�E�P�M�Q�U R�EPj�M$Q���t#�U�R�E�P�M�Q�U�R�EP�MQ�Sn�����EȋU�R�hO�����E�P�\O�����EȋM�3��JV����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�E��M�M��U��U�E����E��}� t�M����t�E����E��֋E+E�����]������������������������U����EP�M���?���M$Q�U R�EP�MQ�UR�EP�MQ�M�� ���P�D����� �E��M���O���E���]��������������������������������U����E�    �E��   �E�;E�A�E�E��+����E��M��U+�x+�U�u�E���}� }�E����E��	�M����M�뷃����]�����������������������������U����E�X$�E�    �E��   �E�;E�W�E�E��+����E�jU�M��U���P�MQ�8�����E�}� u�U��E��D���}� }�M����M��	�U����U�롃����]������������������������������������������������U��Q�   k�����3���U�t#j j j �EP�MQ�UR�EP�MQ�UR�U��'�EP�MQ�UR�EP�MQ�UR�B����P����]��������������������������������������U����} t�}   t	�}   u3��   �} u�} �} }3��   �EP�O�����E��}� }3��i�M���|+�U�jU�E�P�Cp�����E�} ~?�M�;M|3��9j h�   h @hd@h�@�U�R�EP�MQ�rz����P�>�����E����]�������������������������������������������������������������U��Q�} u3��,�EP�1u�����E��}� |	�}��   r3��
�M���x+��]�������������������U��j j �EP�|�]� �����������U����E�    �   k�����3���U�tj �EP�MQ�UR�U��%�E�|�jh����E��|�    �E���]�������������������������������U��Q�   k�����3���U�tj �EP�MQ�UR�EP�MQ�UR�U��'�EP�MQ�UR�EP�MQ�UR�@����P����]��������������������������U��Q�   k�����3���U�t�EP�MQ�UR�EP�U���MQ�UR�EP�MQ�?����P����]����������������������������U��Q�   k�����3���U�t�EP�MQ�UR�EP�MQ�UR�U��'�EP�MQ�UR�EP�MQ�UR�,?����P����]����������������������������U��Q�   k�����3���U�t�EP�MQ�U���UR�EP��P��V������]����������������������������U��Q�   k�����3���U�t	�EP�U��j�MQ�r>����P����]������������������U��Q�   k�����3���U�t#j j j �EP�MQ�UR�EP�MQ�UR�U��'�EP�MQ�UR�EP�MQ�UR��=����P����]��������������������������������������U����E�    �} ��   �E���A|�U���Z�M��� �U��	�E��M�f�U�f�U��E���A|�U���Z�M��� �U��	�E��M�f�U�f�U��E���E�M���M�U���Ut�E���t�M��U�;��a����E��M�+��E�E��]�������������������������������������������������������U����} ~�EP�MQ��j�����E�} ~�UR�EP��j�����E�} t�} u4�M+Mu	�E�   ��U+Uy	�E�   ��E�   �E��E��E�� �MQ�UR�EP�MQ�UR�EP�Vd������]�����������������������������������������������������U��} ~�EP�MQ�,j�����E�UR�EP�MQ�UR�EP�MQ�(����]�������������������U��j�h��h�Ld�    P��$SVW���1E�3�P�E�d�    �e��E� �E�  �E�EЍE�E��E�    �E�Pjj h�m@�8��E� 3Ɂ8�m@����Ëe��E������E�M�d�    Y_^[��]����������������������������������������U��j�h��h�Ld�    P��$SVW���1E�3�P�E�d�    �e��E� �E�  �E�EЋE�EԋE�E؍E�E܋E�E��E�    �E�Pjj h�m@�8��E� 3Ɂ8�m@����Ëe��E������E�M�d�    Y_^[��]������������������������������������������������������U���H  ���3ŉE��EW�=`��������E����������2  S��Vh   j h`F�Ӌ���u"����W��   VVh`F�Ӌ�����   h|FV���ȉ������   ����������   ����   �C�s h�F�u��$h�FPh GVh,Gh@G������h�GP�ыC��$PV�E�P�E�P�  ��8�E�h�GPh�G�E�P������h�GP�  ��������P���������PjW�������  ��(^[_�M�3��I����]�h�FjW��������  ��^[�M�3�_��H����]�����������������������������������������������������������������������������������������������������������U��E��w#��P��� A���t.RPQ�u�7  ��]Ë4A�   RP�   Q�u�  ��]�����������������������������������U���  ���3ŉE��E�������X�������S�]�����   �; ��   S�  ��-��=   ��   3����$    ���PA�@��������u�VW��C��u�������+�O�GG��u��˺lA���˃���B��u�������+�O�GG��u��ʍ��������ʃ��_^��0FPj�������������  ���M�3�[�G����]�����������������������������������������������������������������U��Q�U�MSVW�}3�+׉U�E�M���r�   ;�s%�:��Ph\�Q����M����UF���G�ǋE_� �E�p� ^[��]�����������������������������������������U��U�@��u�+�H]�������������U���<  ���3ŉE��ES�]V�uWV������������ǅ����    �I��������uV�,A����������j j j�S�j h��  ��=   s#P������Pj�������j h��  �Ӎ�������u�Eh  �~�������t$������SV�4�8AP�"��������  2��������� u����   ��t� ����   h  ������P������Ph  ������P�F�P�Ue������t*S������������h�EP������������P�u���   �������j j h
  Pj���������EPj h��  �Ӆ�t������j j h
  ��������EPj�������Pj h��  �Ӆ�t������������������hFV������W�u����������u̋M�_^3�[�"D����]����������������������������������������������������������������������������������������������������������������������������������U���  ���3ŉE��\�������S�]�����   ����   S�7�����:��=   w3����    ���A�@��������u�VW��C��u�������+�O�GG��u��˺�A���˃���B��u�������+�O�GG��u��ʍ��������ʃ��_^���GP�Ej������P�������M�3�[�B����]������������������������������������������������������������������̡������������̡�������������U��E��w	��H]�3�]��������̸   �����������U�졄��M������    ]��������������������U�졈��M������    ]��������������������U��U��w��P��M��P�]Ã��]��������������U��&]�������U�츠%]�������u�U��� PRSVWh�Hh�aj7h�Ij��"������u�_^[ZX��]�������������������������U��j�s^������tj�d^������u#�=��uh�   �L����h�   ��K����]����������������������������U��Q�E�    �	�E����E��}�s�M��U;�(Ju�E���,J���3���]������������������U���   ���3ŉE��EP�M+���������������� �  ǅ����    �}�   t\�}�   tS�}tM������Qhpjj j j j�3!���������������� t������t��ǅ����   �
ǅ����   ������ �  j�]������tj�	]��������   �=����   j��������������� ��   ���������   ǅ ���    ��� ������� ����� ����  s4�� ����� ����������J������� ����������P��u�뱺   i��  �������������  s���^��������Ƅ��� j ������R�����P� J����P�����Q������R����  �}�   ��  �   k���������������������  +����������������j h  h�Uh Vh Vh�Vh  h���f����P�>*�����   i�  3ɋ����f�h  �����Pj �(��u:j h  h�Uh Vh0Wh�������Q�����R�Bf����P��)����������P�H��������<vk�����Q�H�����������DB�������j h#  h�Uh Vh�Wjht�������+������������+�R������P�<5����P�S)����j h&  h�Uh VhXXh��h  h���af����P�)����j h'  h�Uh Vh�X������Qh  h���)f����P��(����h  h��h���=�����M�3��<����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE��}��  �E��h�����|�����x���ǅd���    ǅl����   ��l���R��x���P�MQ�UR�EP�df������p�����p��� ��   ����zt�/  j j �MQ�UR�EP�)f������l�����l��� u�  j^h�Yjj��l���Q�4������x�����x��� u��   ǅd���   ��l���R��x���P�MQ�UR�EP�e������p�����p��� u�   jih�Yjj��p���Q�24������h������h����8 u�fj jlh�Yh4Zh`Z��p�����Q��x���R��p���P��h����R�{g����P�6&������d��� tj��x���P��)����3��6  ��d��� tj��x���Q��)��������  �  �}��   �U��t�����t����     j j �MQ�UR��������`�����`��� u�\h�   h�Yjj��`���P�/3������t������t����: u�*��`���P��t����R�EP�MQ�y������u�3��oj��t����P�)������t����    ����K�F�} u@ǅ\���    j��\���R�E    P�MQ�������u�����U��\����3������M�3���8����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E���]����U����E�    �} t	�E�   ��E�    �E�E��}� u&h\hpjj hJ  h[j��������u̃}� u3�)_���    j hJ  h[h,\h\�tW�����   �R  �} t	�E�   ��E�    �U�U�}� u&hl\hpjj hK  h[j�S������u̃}� u3�^���    j hK  h[h,\hl\��V�����   ��   �����u����u�E�   �M�    j j j��URj �E�P��E��}� u��P�����3��|h\  h�\j�M���Q������U��E�8 u3��Q�M�Q�U�Pj��MQj �U�R���u,��P�/����j�E�Q��%�����U�    3���   ��]�����������������������������������������������������������������������������������������������������������������������������U����E�    �} t	�E�   ��E�    �E�E��}� u&h�\hpjj h�  h[j�t������u̃}� u3��\���    j h�  h[h�\h�\�U�����   �X  �} t	�E�   ��E�    �U�U�}� u&h]hpjj h�  h[j��������u̃}� u3�H\���    j h�  h[h�\h]�T�����   ��   �%����u����u�E�   �M�    j j j j j��URj �E�P��E��}� u��P�)����3��~h�  h�\j�M�Q�Q�����U��E�8 u3��Uj j �M�Q�U�Pj��MQj �U�R���u,��P������j�E�Q�#�����U�    3���   ��]���������������������������������������������������������������������������������������������������������������������������������������U����E�Ph�Zj �,��th [�M�Q���E��}� t�UR�U���]�������������������U��EP�84�����MQ��]����������������������U������P��E��$��M��	�U����U��}� t�E��8 tj�M��R�2"������j�$�P� "�����$�    � ��M��	�U����U��}� t�E��8 tj�M��R��!������j� �P��!����� �    j��Q�!����j��R�!������    ��    �}��t�=�� tj�E�P�u!����j������   k� ��,� t+j�   k� ��,�R�>!�����   k� ǁ,�    �   �� ��,� t+j�   �� ��,�Q�!�����   �� ǂ,�    �|������Iu'�=|�X�tj�|�R�� �����|�X���]������������������������������������������������������������������������������������������������������������������������������U���zQ���EP�i;����h�   ���]�����������������U��jjj �B  ��]��������������U��jj j �"  ��]��������������U��Q�=�� th����Q������t�EP������B��h�Xh�V�*�����E��}� t�E��Gh'q�7����h�Uh P��  ���=t� tht��lQ������tj jj �t�3���]������������������������������������������������������U��j j�EP�0  ��]������������U��j j j �  ��]��������������U����} t	�E�   ��E�    �E��E��}� u&h��hpjj h%  h[j��������u̃}� u3� V���    j h%  h[h�[h���kN�����   �   �=(� t	�E�   ��E�    �U�U��}� u&h�[hpjj h)  h[j�G������u̃}� u0�U���    j h)  h[h�[h�[��M�����   ��M�(��3���]������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u&h��hpjj h  h[j�k������u̃}� u3��T���    j h  h[h�[h���M�����   �   �=,� t	�E�   ��E�    �U�U��}� u&h�[hpjj h  h[j��������u̃}� u0�<T���    j h  h[h�[h�[�L�����   ��M�,��3���]������������������������������������������������������������������������U��Qj ��E��E�P�)�����M�Q�$�����U�R�������E�P�6�����M�Q�@�����U�R�U�����(G����]���������������������������������U��E;Es�M�9 t�U��ЋM���M��]����������U��Q�E�    �E;Es#�}� u�M�9 t
�U��ЉE��M���M�ՋE���]��������������������U��j�@����]������������������U��j�yE����]������������������U��j�hИh�Ld�    P���SVW���1E�3�P�E�d�    �����E�    �=0��N  ��   �E���} �  ���Q��E��}� ��   ���R��E��E�    �E��E؋M�Mк   ����   �E�    �E�    �E���E�M�;M�rj ��U�9u�ދE�;E�s�k�M�R��E�j ��M��Ű��R��Eܡ��P��EԋM�;M�u�U�;U�t�E܉E؋M؉M��UԉUЋEЉE��N���h�\h�Y�������h�^h�]��������} uj���/������ t
�3(����B���E������   ��} t�#)��Ã} t��0�   �)���MQ�4�����M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������U��j j �EP������]������������U����E�8�t%�M��E��M��U�EB3E��E��M��*(���M�Q�E��M��U�EB3E��E��M��(����]������������������������������������U���0�E� �E�   �E���E��M����M�U��B3���E�M�Q�U�R�A������E�H��f�  �U�UЋE�EԋM��UЉQ�E��H�M���U܉U��}����   kE��M�T�U�E�H�M�U��E܃}� ��   �U�M��1���E��E��}� }�E�    �   �   �}� ��   �M�9csm�u)�=� t h���H������tj�UR�����M����U�I���E��H;M�th���U�R�M����U�����E��M܉H�U�R�E�P�)������U�M�I��$�������&�U��z�th���E�P�M���������/���E��M���t�U�R�E�P��������E؋�]�����������������������������������������������������������������������������������������������������������������������������U��   ]�������U���h�    ]������������������U���E%�  ���ȋU�����P���E�$������]�����������������U����E��������Dz���]��E�    ��   �E%�  ��   �M����u
�} ��   �E�������]����Au	�E�   ��E�    �U��U��E��u/�M��M�U��   �t	�E���E�M��M�U����U����E%��  f�E�}� t�M�� �  f�Mj ���E�$������]��.j ���E�$�������]��U���  ����-�  �E��M�U���E��]����������������������������������������������������������������������������������U��Q�E%�  ��f�E��M����  f�M��E���]�����������������������U����E�]��E%�  �M���f�E��E���]�������������������������U����E�]�E�  �E��M���  �U����f�M��E��]�����������������������������U��}  �u�} u�   �X�}  ��u�} u�   �B�E%�  =�  u�   �+�M���  ���  u�U����u�} t�   �3�]������������������������������U��Q�E�� t	�E�   �K�M��t	�E�   �:�U��t	�E�   �)�E��t	�E�   ��M��t	�E�   ��E�    �E���]��������������������������S�܃������U�k�l$���   ���3ŉE��C P�KQ�SR��������u)�E�����E��KQ�SR�CP�KQ�S R�E�P�	�����KQ�������|����=P� u>��|��� t5�S R���C�$�����$���C�$�CP��|���Q�D����$�%���|���R�/����h��  �C P�"2�����C�M�3�� !����]��[�����������������������������������������������������������������������������S�܃������U�k�l$���   ���3ŉE��C(P�K Q�SR�������u;�E����E��M������M��C�]��S R�CP�KQ�SR�C(P�M�Q������SR�c������|����=P� u?��|��� t6�C(P���C �$���C�$���C�$�KQ��|���R������$�%���|���P�=.����h��  �K(Q��0�����C �M�3������]��[��������������������������������������������������������������������������U��Q�E�    �	�E����E��}�}�M��͠�;Uu�E��Ť����3���]������������������U���H�E���E��M��t �U��tj��8�����E�����E��  �M��t �U��tj��8�����E�����E��s  �M���   �U���  j�8�����E%   �E�}�   w�}�   tW�}� t �}�   tv��   �}�   ��   �   �M�������z�p��]���p����]ЋU�E���   �E�������z�p��]��������]ȋM�E���Z�U�������z����]���p����]��E�E���,�M�������z����]��������]��U�E���E�����E��G  �M���;  �U���/  �E�    �E��t�E�   �M���������D��   �U�R�E��� �$�K�����]؋M��   �M��}�����}�E���s�]��E�   �   ���]�����Au	�E�   ��E�    �U�U��Eރ�f�E��Mރ�f�M��	�U����U��}����}:�E؃�t�}� u�E�   �M���M؋U܃�t�E�   ��E؋M���M�봃}� t�E����]؋U�E����E�   �}� t
j�Z6�����E�����E��M��t�U�� tj �76�����E����E��}� t	�E�    ��E�   �E��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��=P� u0�EP���E�$�����$���E�$�MQj�����$�!��B��� !   h��  �UR��+�����E]������������������������������������U����E�E�]��=P� u1�EP���E��$���E�$���E�$�MQj�{
����$�!���A��� !   h��  �UR�]+�����E���]�������������������������������������U��j �EP�MQ�UR�EP�MQ�UR�z,����]����������U���,�E�  ��E�@    �M�A    �U�B    �E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U��t�E��  ��E�H���U�J�E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U���t	�E�    ��E�   �M�����U�B�����M�A�U���t	�E�    ��E�   �M�����U�B�����M�A�U���t	�E�    ��E�   �M������U�B�����M�A�U���t	�E�    ��E�   �M܃���U�B�����M�A�U��� t	�E�    ��E�   �M؃��U�B�����M�A��,���E��U���t�E�H���U�J�E���t�M�Q���E�P�M���t�U�B���M�A�U���t�E�H���U�J�E��� t�M�Q���E�P�M���   �U�}�   w�}�   t+�}� tI�}�   t.�K�}�   t�@�E����U�
�1�E�������U�
��E�������U�
��E�����U�
�E���   �M�t5�}�   t�}�   t�1�U����M��"�U������M���U������M��U���  ���E��� ��ʋU�
�}  tT�E�H ���U�J �E�H ���U�J �E�M��X�U�B`���M�A`�U�B`���M�A`�U�E� �ZP�X�M�Q ���E�P �M�Q �����E�P �M�U��Y�E�H`���U�J`�E�H`�����U�J`�E�M��XP�����URjj �E�P�8�M�Q����t�E�����U�
�E�H����t�U�����M��U�B����t�M�����E��M�Q���t�E����U�
�E�H��t�U���ߋM��U����Eԃ}�w[�M��$��/�U�%����   �M��;�U�%����   �M��%�U�%����   �M���U�%�����M��U������E�t�}�t �}�t2�@�M���������   �E��(�M���������   �E���M��������E��}  t�M�U�BP���E�M�AP���]ÐT/>/(//����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�EP�MQ�UR�EP�MQ�UR�j%����]����������U��Q�E�E��}�t�}�~ �}�~��V:��� !   ��I:��� "   ��]�����������������������U��� �EP�!������E�}� t^�M�M��U�U�E�E�M�M��U�U�E �E��M$�M�h��  �U(R�L#�����E�P�������u�MQ� �����E��"� h��  �U(R�#�����EP�i �����E ��]����������������������������������������������������U��Q�=@�|�*���E��E���?�E�������E�    �E���]��������������U����=@�|8�����E��E#E�M��#M���E��U������U��U��E�P��������E�    �E���]����������������������������U��Q�=@�|�]��e���U���]��������������������U��Q�=@�|�]���E�    �E���]����������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �e�=@���   �E��@tp�=к tg�E�    �U�E������Q�M���E�}�  �t�}�  �t	�E�    ��E�   �E�Ëe��к    �M�ΈM�U�E�������U�⿉U�U�M�d�    Y_^[��]����������������������������������������������������������U��Q����E��E��?E��E��M�Q���������]�������������������������U��Q�=@�|�����E��E���?�E���E�    �E���]�������������������U��Q�}����E���]����������������U�����}��E#E�M��U��#��f�E��m��E���]���������������������U����E��t
�-���]���M��t����-���]������U��t
�-ĺ�]���E��t	�������؛�M�� t���]����]����������������������������U��Q��}��E���]�����������������U���0���3ŉE�SV�@�    �ܺ���ܺj
�v�����[  �E�    �E�    �E�    �@�   �ܺ���ܺ�u�3�3����^�N�V�   k� �L��Mк   �� �D�5Genu�   k��L���ineI��   ��L���ntel�u	�E�   ��E�    �UԈUߍu�   3����^�N�V�   k��   k� �L��L�   ��   �� �L��L�   k� �L��M��U߅�to�E�%�?�=� tS�M؁��?���` tB�U؁��?���p t1�E�%�?�=P t"�M؁��?���` t�U؁��?���p u�D����D��}�|O�u�   3����^�N�V�   �� �   ��D��D�   �� �T���   t�D����D��   �� �T���   ��   �@�   �ܺ���ܺ�   �� �T���   tV�   �� �L���   tB�@�   �ܺ���ܺ�   ���L��� t�@�   �ܺ�� �ܺ3�^[�M�3��|����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̅�uf���fn�f`�fa�fp� SQ�ك���ux�ڃ���t0ffAfA fA0fA@fAPfA`fAp���   KuЅ�t7����t��I f�IKu���t����t
f~�IJu���t�AKu�X[��ۃ�+�R�Ӄ�t�AJu���t
f~�IKu�Z�^�����������������������������������������������������������U���0�} t�} v	�E�   ��E�    �E�E��}� u#h^hpjj jhx^j��������u̃}� u0�1���    j jhx^h�^h^�[)�����   �k  �} ��   �U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U�E�Ph�   �M��Q�-�����} t	�E�   ��E�    �U�U�}� u#h�^hpjj jhx^j���������u̃}� u0�30���    j jhx^h�^h�^�(�����   �  �M�M��U�U��E��M���E���MЋU����U��E���E�}� t�M����M�t�ȃ}� ��   �U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U��E�Ph�   �M��Q������ _��t3�t	�E�   ��E�    �M܉M؃}� u#hP_hpjj jhx^j��������u̃}� u-�/��� "   j jhx^h�^hP_�\'�����"   �o�}�tg�}���t^�E+E���;EsP�M+M����U+�9h�s
�h��E���M+M����U+щUԋE�Ph�   �M+M��U�D
P�#����3���]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u#h�hpjj j)h�_j���������u̃}� u+�S-���    j j)h�_h�_h��%���������U�B��]�������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u�����     �,��� 	   �����  �} |�E;\�s	�E�   ��E�    �M��M܃}� u#h`hpjj j.h�`j���������u̃}� u9�*����     �8,��� 	   j j.h�`h�`h`�$��������9  �E���M������P��D
��t	�E�   ��E�    �M؉Mԃ}� u#h�`hpjj j/h�`j�P�������u̃}� u9�����     �+��� 	   j j/h�`h�`h�`��#��������   �EP�E0�����E�    �M���U������P��L��t�UR������E��9�(+��� 	   �E�����3�u#h(ahpjj j9h�`j��������u��E������   ��UR�+�����ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������U��QV�EP���������tn�}u�   k� ��P����   ��u�}u1�   k� ��P��QD��tj�H�������j�<�����;�t�EP�,�����P����t	�E�    �	���E��MQ�}������U���E������P��D �}� t�U�R����������3�^��]����������������������������������������������������������������������U��} u#h�ahpjj j.h bj�}�������u̋M�Q��   tK�E�H��t@j�U�BP��������M�Q�������E�P�M�    �U�B    �E�@    ]������������������������������������������U��j�h0�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u�(��� 	   �����  �} |�E;\�s	�E�   ��E�    �M��M܃}� u#hhbhpjj j,h�bj�Y�������u̃}� u.�'��� 	   j j,h�bhPchhb����������X  �E���M������P��D
��t	�E�   ��E�    �M؉Mԃ}� u#hdchpjj j-h�bj���������u̃}� u.�'��� 	   j j-h�bhPchdc�i���������   �EP��+�����E�    �M���U������P��L��t;�UR�/�����P����u���E���E�    �}� u�C�p����M��&��� 	   �E�����3�u#h(ahpjj jEh�bj���������u��E������   ��MQ������ËE�M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������U��j�hP�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u�.����     �<%��� 	   �����  �} |�E;\�s	�E�   ��E�    �M��M܃}� u#h`hpjj jBh�cj�~�������u̃}� u9�����     ��$��� 	   j jBh�chdh`���������L  �E���M������P��D
��t	�E�   ��E�    �M؉Mԃ}� u#h�`hpjj jCh�cj���������u̃}� u9�����     �*$��� 	   j jCh�chdh�`�x��������   �EP��(�����E�    �M���U������P��L��t�UR�EP�MQ��������E��D�#��� 	   �����     �E�����3�u#h(ahpjj jNh�cj��������u��E������   ��MQ������ËE�M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������U�츔<  �")�����3ŉE�ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    �} u3��C  �} tǅ|���   �
ǅ|���    ��|��������������� u#hdhpjj jlh�cj��������u̃����� u9������     ��!���    j jlh�ch<dhd�4��������  �U���E������P��T$������������������t����������   �U��uǅ����   �
ǅ����    ��������x�����x��� u#h`dhpjj jth�cj���������u̃�x��� u9� ����     �!���    j jth�ch<dh`d�\���������  �U���E������P��T�� tjj j �EP������MQ���������   �U���E������P��T��   tt�O����p�����p����Hl�   �⃼�    uǅ����   �
ǅ����    ��������������l���Q�U���E������P��R�������������� �  ������ t����������  ����t���3�f������ǅ����    ǅ����    �U������������+E;E��  ǅ����    ���������  ���������
uǅ����   �
ǅ����    �������������U���E������P��|8 ��   �U���E������P��T4R�R"������u&h�dhpjj h�   h�cj��������u̋M���U������P��   k� �T4�T��   �� ��������T�E���M������P��D
8    j�E�P������Q�I��������u�{  ��   �������P�!��������   ������+M�U+у�v3j������P������Q����������u�'  ���������������T�E���M������P�������� �D
4�M���U������P��D8   ����������������  �"j������R������P�l��������u�  ���������������e��������t��������uM������f�f��������������
uǅ����   �
ǅ����    �����������������������������������P  j j j�M�Qj������Rj ��t���P������������� u��  �sj ������Q������R�E�P�M���U������P��Q����t*������+U�����������������;�����}�  ����������n  ������ ��   ǅ����   �   k� �D�j ������P������Q�U�R�E���M������P��
P����t3������;�����}��   ���������������������������������������   ��   ��������t����������   ������P�������������;�u������������������������p������ tbǅ����   �   f������������R��������������;�u ���������������������������������������D����7  �M���U������P��L��   ��  ǅ����    ���������[  ǅ����    ǅ����    �E������������+M;M�'  ������������������������+�=�  ��   ������+U;Usr�����������������������������������
u'���������������������������������������������������������������g���j ������Q������������+�R������Q�U���E������P��R����t,�����������������������������+�9�����}�����������������A  ���������[  �M������ǅ����    ������+U;U�1  ������������������������+ʁ��  ��   ������+E;Es{������f�f����������������������������
u,���������������   ������f���������������������f������f����������������]���j ������P������������+�Q������P�M���U������P��Q����t,�����������������������������+�9�����}�����������������  �U������ǅ����    �E������������+M;M��  ǅ����    ��H�����������������H���+�=�  sz������+U;Usl������f�f����������������������������
u�   ������f�
��������������������f������f����������������q���j j hU  ������Q��������H���++���P��H���Pj h��  ������������� u���������   �   ǅ����    j ������Q������+�����R������������Q�U���E������P��R����t���������������������������������;������������;�����~�������+E�������F����Yj ������Q�UR�EP�M���U������P��Q����tǅ����    ��������������������������� ��   ������ t9������u���� 	   �q�����������������R�����������\�L�E���M������P��D
��@t�M���u3��+��4���    �����     �����������+������M�3��j�����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���V�E�    �} t	�E�   ��E�    �E��E�}� u#hl�hpjj jmh�dj���������u̃}� u.�;���    j jmh�dh4ehl��	���������  �U�U��E��H��   t�U��B��@t����  �M��Q��t�E��H�� �U��J����  �E��H���U��J�E��H��  u�U�R��������E��M��Q��E��HQ�U��BP�M�Q�{�����P�A������U��B�E��x t	�M��y�u:�U��z t	�E�    ��E�   �E��HM��U��J�E��@    �����   �M��Q��   u�E�P���������t@�M�Q����������t/�U�R������������E�P������������P��E���E���M��Q��   ���   u�E��H��    �U��J�E��x   u#�M��Q��t�E��H��   u
�U��B   �E��H���U��J�E������   �U�E�����U��
�E�^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hp�h�Ld�    P�ĄSVW���1E�3�P�E�d�    j��������E�    h�   hHejj@j �H������E�}� u"�E�����j��E�Ph���������E��G  �   k� �E䉂P��\�    �	�M��@�M�   k� ��P���   9M�su�U��B �E�� �����M��A
�U��B    �E�H$�ဋU�J$�E�H$���U�J$�   k� �U��D
%
�   �� �M��D%
�U��B8    �E��@4 �i�����t���Q���U�����  �}� ��  �E���M܋U����UԋE�E܉E؁}�   }�M܉M���E�   �UĉU��E�   �	�EЃ��EЋ\�;M���   h�   hHejj@j ��������E�}� u�\��U��   �EЋM��P��\��� �\��	�E��@�E�MЋ�P���   9U�sf�E��@ �M�������U��B
�E��@    �M�Q$�​E�P$�   k� �E��D%
�   �� �U��D
%
�E��@8    �M��A4 �|��������E�    ��U����U��Eԃ��EԋM؃��M؋U�;U���   �E؃8���   �M؃9�ty�U����tn�M����u�E؋Q����tS�U����E������P��E�M�U؋��M�UԊ�Aj h�  �M��Q�l������U�B���M�A�G����E�    �	�U����U��}��H  �   k� �U����P��U�E�8�t�M�9��  �U��B��}� u	�E�������}�u	�E�������E������E��E��M�Q���Ẽ}����   �}� t�U�R���Eȃ}� tl�E�M̉�Uȁ��   ��u�E��H��@�U�J��E�%�   ��u�M��Q���E�Pj h�  �M��Q�T������U�B���M�A�5�U��B��@�M�A�U�������=� t�E������B������E��H�ɀ   �U�J�����E������   �j�������3��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    �	�E����E��}�@}y�M��<�P� tg�U���P��E��	�M���@�M��U���P�   9E�s�M��y t�U���R���j�E���P�Q�%������U���P�    �x�����]������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�   ��E�    �E�E��}� u#h�hpjj j0hxej��������u̃}� u.����    j j0hxeh�eh��Y������������F�UR�������E�    �EP�'������E؉U��E������   ��MQ�s�����ËE؋U܋M�d�    Y_^[��]����������������������������������������������������������������������������������U��\  ������3ŉE�V�} u#hl�hpjj jZhxej蘿������u̋M������������R��������������������x }�������A    jj j ������R�W����������������������� |	������ s�������[  ��������������������P��D
$�����������������Q��  u#�������@�������+ȋ�����������  �������������
+H�������������B���  ����������  ��������������������P��|0 �m  �������������
+H�鉍�����������z u�������������g  �2  j ��������������������P��D
,P�L
(Q������R���������������������������������������P�������������������������������;T(u������������������;T,t�������  j ������Ph   ������Q��������������������P��R����u�������r  j ������P������Q������R�$����������������������� |	������ s�������(  ������;�����v�������  �������������������������������������������� ��   ������������9�����ss���������u5������������9�����s�������Q��
u������������������������X���������������������������P���������������+Ћ�3������������0  ��������������������P��L��   tO�������B���������������������������������;s���������
u�����������������'�������Q��   u�����    �������  �����������u3ҋ������t  �������Q���4  �������x uǅ����    �  �������������+B������A��������������������������P��T��   ��  jj j ������P������������������������;�������   ������;�������   �������H������������������B���������������������������;�����s���������
u���������������ċ������H��    t����������������   j ������P������Q������R������������������������� |	������ s��������   ������   w*�������H��t�������B%   uǅ����   ��������Q��������������������������P��D
��t����������������������u�������艅����3ɋ�����+��������������������������������u�������ꉕ����������3�����������^�M�3�������]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} u#hl�hpjj jdh�ej躶������u̋M�M��U�R�
������E��E��H��   u$������ 	   �U��B�� �M��A����X  �-�U��B��@t"������ "   �M��Q�� �E��P����)  �M��Q��tH�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J�����  �E��H���U��J�E��H���U��J�E��@    �E�    �M�M��U��B%  uC�����    �� �9E�t�u����    ���9E�u�E�P�V�������u�M�Q�$������U��B%  ��   �M��U��+By&h`fhpjj h�   h�ej�*�������u̋U��E��
+H�M�U��B���M���U��B���M��A�}� ~�U�R�E��HQ�U�R�k������E��q�}��t!�}��t�E����M������P��M���E���U��B�� t7jj j �M�Q�������E�U�U�#U���u�E��H�� �U��J����O�E��H�U���E�   �E�P�MQ�U�R��������E��E�;E�t�M��Q�� �E��P�����E%�   ��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E������E������}�u!�W����     �e���� 	   ��������  �} |�E;\�s	�E�   ��E�    �M�M��}� u#h`hpjj j@h�fj褲������u̃}� u<�����     ������ 	   j j@h�fh\gh`�<������������`  �E���M������P��D
��t	�E�   ��E�    �M܉M؃}� u#h�`hpjj jAh�fj��������u̃}� u<�?����     �M���� 	   j jAh�fh\gh�`�������������   �EP��������E�    �M���U������P��L��t �UR�EP�MQ�UR�������EЉU��K������ 	   襶���     �E������E�����3�u#h(ahpjj jLh�fj�#�������u��E������   ��UR躮����ËEЋUԋM�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EP�������E��}��u:����� 	   3�u#h(ahpjj jwh�fj���������u̃������s�EP�M�Q�UR�EP�M�Q����u��P苮�����������>�U���E������P��T����E���M������P��T�E�U���]�����������������������������������������������������U����} u#hl�hpjj j.hxgj��������u̋|����|��U�U�j:h�gjh   ��������E��E��M��H�}� t�U��B���M��A�U��B   �%�E��H���U��J�E����M��A�U��B   �E��M��Q��E��@    ��]������������������������������������������������������������U��j�hЙh�Ld�    P���SVW���1E�3�P�E�d�    �E�    j��������E�    �E�   �	�E���E�M�;���   �U䡜�<� t|�M�����H��   t"�U䡜��Q����������t	�U����U��}�|=�E������ R�j�E����R�������E����    �Y����E������   �j������ËE��M�d�    Y_^[��]���������������������������������������������������������������������������U���0�} t�} v	�E�   ��E�    �E�E��}� u#hhhpjj jhx^j般������u̃}� u0������    j jhx^hthhh�+������   �w  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R��������} t	�E�   ��E�    �E�E�}� u#h�^hpjj jhx^j誫������u̃}� u0������    j jhx^hthh�^�M������   �  �U�U��E�E��M��Uf�f��M���UЋE����E��M���M�}� t�U����U�t�ƃ}� ��   3��Mf��}�tJ�}���tA�}v;�U��9h�s
�h��E��	�M���M��U���Rh�   �E��P�������� _��t3�t	�E�   ��E�    �E܉E؃}� u#hP_hpjj jhx^j耪������u̃}� u-������ "   j jhx^hthhP_�#������"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9h�s�h��U���E+E����M+ȉMԋU���Rh�   �E+E��M�TAR�������3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�E��M�Q�UR�EP�MQ��������]�����������U��Q�E�E��M�Q�UR襭������]�������������������U��Q�E�E��M�Q�UR�EP��������]���������������U��Q�E�E��M�Q�UR��������]�������������������U��Q�E�E��M�Q�UR�EP���������]���������������U��Q�E�E��M�Qj �UR�EP�MQ�UR��������]���������������������U��Q�E�E��M�Q�UR�EP�MQ�UR�EP�˲������]�������������������U���L�E�    3��E��E��E��EĉEȉẺEЍM��M��} t	�E�   ��E�    �U��U�}� u&h��hpjj h�   h�hj�'�������u̃}� u1�|����    j h�   h�hh�hh�������������o  �} t	�E�   ��E�    �M��M�}� u&hX�hpjj h�   h�hj訦������u̃}� u1������    j h�   h�hh�hhX��H����������   �E�E܋M��AB   �U��E�B�M��U��E��@����M�Qj �UR�E�P�e������E��} u�E��   �M��Q���U�E��M�H�}� |"�U���  3Ɂ��   �M؋U�����M����U�Rj � ������E؋E��H���M�U��E�B�}� |!�M��� 3�%�   �EԋM�����E����M�Qj ��������EԋE���]�����������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�E��M�Qj �UR�EP�MQ胮������]�������������������������U��Q�E�E��M�Q�UR�EP�MQ�UR�A�������]�����������������������U��Q�E�E��M�Q�UR�EP�MQ�UR蟫������]�����������������������U��Q�E�E��M�Qj �UR�EP�MQ�a�������]�������������������������U��������d]����U�졌�P�]����������������U���������`]����U��E����M����U����E���]����������U��j�h0�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    j �%������E�    �} u�E����E��Q��E��E�   ��E����U��P��E��E�   �}� t�}�tj ��M���E������   �j ������Ã}� u3���}�t
�U�R�U���   �M�d�    Y_^[��]� ��������������������������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�    �E�    �E�    �E�    �E�EԋMԃ��Mԃ}���   �U������$�l��E���M��U��E؃��E��  �E���M��U��E؃��E���   �E���M��U��E؃��E���   �E���M��U��E؃��E��   �����E܃}� u�����  �M܋Q\R�EP��  �����E�M��U��   �}3�t	�E�   ��E�    �M̉Mȃ}� u&h<ihpjj h�  h�ij轠������u̃}� u1�����    j h�  h�ih�ih<i�]���������5  �E�P��E��}�u3��  �}� uj�c����}� t
j �C������E�    �}t�}t�}u,�M܋Q`�UċE��@`    �}u�M܋Qd�U��E��@d�   �}u:�H��M��	�UЃ��UСH�L�9E�}kM��U܋B\�D    ���j ��M��E������   ��}� t
j �������Ã}u�U܋BdPj�U����
�MQ�U����}t�}t�}u�U܋EĉB`�}u	�M܋U��Qd3��M�d�    Y_^[��]Ë��h�.�K���� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�E��M��Q;Ut�E����E�k@�M9M�s��k@�U9U�s�E��H;Mu�E���3���]���������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�    �}t�}u�R  �}t�}t�}t�}t
�}�F  j �;������E�    �}t�}u=�=�� u4jh0�����u���   ������G����0�E�   �E�E؋M؃��M؃}���   �U���X��$�D����Q��E܃}t�UR�����r���P��E܃}t�MQ�����L���R��E܃}t�EP�����%���Q��E܃}t�UR�����E������   �j �i�����Ã}� t��   ��   �}t�}t�}t��   �U����E��}� u��   �E��x\��uLhZ  hij�D�Q������E̋U��ẺB\�}� t�D�Qh���U��B\P�Ӥ������h�M��Q\R�EP�@������E�}� u�J�M�Q�U܃}t3�E�H;Mu(�U�E�B�M���M�k@��E�P\9U�r��͋E��   �M�MԋUԃ��Uԃ}�w�E���x��$�p�����}3�t	�E�   ��E�    �EȉEă}� u&h<ihpjj h�  h�ij谚������u̃}� u.�����    j h�  h�ih�ih<i�P�������������M�d�    Y_^[��]Ë�܈)�P��u� �I ����     �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���`���3ŉE��E�    j ��E��E�    �E�    �d����E��E�    �=�� ��   h   j hj���E�}� u����Wuj j hj���E�}� u3��q  h$j�E�P���E�}� u3��R  �M�Q����h4j�U�R��P����hHj�E�P��P����h`j�M�Q���E�U�R�����=�� th�j�E�P��P����� ��t �} t
�MQ���}� t
�   �  �}� ��   ���R��E��E�    �E��E��M�M��U�U��E�E�3ɉM��}� u3��S  j j �U�Rh�*j j ���E؃}� u3��,  j j��E�P����u�E��  3��  ���;M�th���;U�t]���P��Eԋ��Q��E��}� t8�}� t2�UԉE܃}� t�U�Rj�E�Pj�M�Q�U���t�U���u�E�   �}� t�E    �E�W���;M�t���R��E��}� t�U��E�}� t*���;E�t ���Q��EЃ}� t
�U�R�UЉE䡨�P��Eȃ}� t�MQ�UR�EP�M�Q�U���3��M�3�������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�E��M��QR�E��HQ�U��BPj �M���ҋM��A3���]� ��������������������������U���]�����������U��X�]�������U����} |�}}	�E�   ��E�    �E��E��}� u*h�jhpjj h�   h kj腔������u茏���}� u0������    j h�   h kh�lh�j�!�����������c�}�u�U��8��Q�E��8��M�}�uj����U��8��'�}�uj����M��8���U�E��8��E��]����������������������������������������������������������������������������U��Q�X��E��M�X��E���]���������������������U����} |�}}	�E�   ��E�    �E��E��}� u'h�jhpjj jsh kj��������u�����}� u.�i����    j jsh kh`kh�j����������   �}�t�U���t	�E�    ��E�   �E�E��}� u'h�khpjj jxh kj蓒������u蚍���}� u+������    j jxh kh`kh�k�2���������/�}�u�U��,���E��,��M�U�E��,��E��]�����������������������������������������������������������������������������������U��j�hP�h�Ld�    P���LP  �������1E�3ŉE�SVWP�E�d�    ǅܯ��    ǅ���    ƅ���� h�  j ������P�u�����ƅ���� h�  j ������Q�X�����3�f�����h�  j �����P�9�����ƅ���� h�  j ������Q�������} |�}|����t  �E�    �}��   �D��   ��@����   j h  h kh�lh�lj
h   ������Q�UR������P�s�����hPm���} t�E�������
ǅ�����m������Q��h�m��������R��h�G���M���ǅܯ�������  �} ��   ǅ̯��    �z���� �������m����     �M Q�URh�  h   ������P��������̯����̯�� }*j h-  h kh�lh��j"j�����Q�	����� �������������̯�� }8j h0  h kh�lh�mhXnh   ������P������P�5������}uV�} tǅ����\o�
ǅ����toj h5  h kh�lh�n������Qh   ������R������P�ٙ����j h7  h kh�lh�o������Ph   ������Q�������P蟙�����}u�U��,���t8j h<  h kh�lh phXph   ������Q������P�R�����j h=  h kh�lh`ph�Gh   ������R�Y�����P�������} ��   ǅЯ��    ����� �������~����     ������Q�UR�EPh�ph�  h   ������Q�a�������Я����Я�� }*j hD  h kh�lh��j"j�����R������ �������������Я�� }8j hG  h kh�lh�phXnh   ������R������P�:������:j hK  h kh�lh�q������Ph   ������Q�������P�������ǅ����    ǅȯ��    j�������Rh   �����P������Q�6�������ȯ��j hP  h kh�lh�qj"j��ȯ��R������ ��ȯ�� t8j hR  h kh�lh�rh�sh   �����P�������P�V������=T� u�=D� �#  ǅԯ��    ǅد��    j�@������E�   �T���ԯ�����ԯ���B��ԯ����ԯ�� tHǅ����    ������Q������R�EP��ԯ���Q�҃���tǅ���   ��������ܯ���렃���� un�D���د�����د���B��د����د�� tHǅį��    ��į��Q�����R�EP��د���Q�҃���tǅ���   ��į����ܯ�����E�    �   �j������Ã���� ��  �=X� t?ǅ����    ������Q������R�EP�X�����tǅ���   ��������ܯ������� �4  �U��,���t>�M�<�8��t1j ������R������P�Ѵ����P������Q�U��8�P���M��,���t������P���M��,�����   �   k� ������������   s�����������Ƅ���� �} t9j h�  h kh�lh�lj
h   ������P�MQ�c�����P�є�����} t�������������
ǅ����    ������P�MQ������R�EP�MQ�UR�o�������ܯ���E������   ��}u�D������Ë�ܯ���M�d�    Y_^[�M�3��6�����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���T�  �������1E�3ŉE�SVWP�E�d�    ǅ���    ǅ���    3�f������h�  j ������Q������3�f�����h�  j �����P�ĭ����ƅ���� h�  j ������Q觭����3�f�����h�  j �����P舭�����} |�}|����v  �E�    �}��   �D��   ��B����   j h�  h khth@tj
h   ������P�MQ������P�ߐ����h�t���} t�U������
ǅ����t�����P��h u��������Q��h4u��蹀��ǅ��������  �} ��   �����������������     �E P�MQh�  h   �����R����������������� }*j h  h khth��j"j����� P������ �~�������������� }8j h
  h khth8uh��h   �����R������P諏�����}uV�} tǅ����v�
ǅ����vj h  h khth�u�����Ph   ������Q������P�O�����j h  h khth w�����Rh   ������P�Y�����P�������}u�M��,���t8j h  h khth�wh�wh   ������P������P�Ȏ����j h  h khth�wh4uh   ������Q�������P萎�����} ��   ǅ���    ����������������     ������P�MQ�URhHxh   h   �����P�)��������������� }*j h   h khth��j"j�����Q脀���� ��������������� }8j h"  h khth��h��h   �����P������P谍�����:j h&  h khthhx������Qh   �����R�������P�t�����ǅ���    j h,  h khth�xj"jj������Ph   ������Qj �B�����P����� ���������� t8j h.  h khth�yhpzh   ������R������P�������=T� u�=D� �!  ǅ���    ǅ���    j�˂�����E�   �T�������������Q���������� tHǅ���    �����P������Q�UR������H�у���t����������ǅ���   �렃���� um�D�������������Q���������� tHǅ���    �����P�����Q�UR������H�у���t����������ǅ���   ���E�    �   �j�"�����Ã���� ��  �=X� t?ǅ���    �����P������Q�UR�X�����t����������ǅ���   ����� �W  �M��,����[  �E�<�8���J  �M��8�R������������t�Jj �����P�����Q輩����P�����R�E��8�Q����t��   ����t��   ǅ���    j h�  h khth�zj"jj������Rh   �����P�����Q聜����P��|���� ���������� t>�����Pt5j �����R�����P�	�������P�����Q�U��8�P���@����� v������������j �����R�����P�����Q�U��8�P���M��,���t�����P���M��,�����   �   k� ����������    s�腽��3ҋ����f�������} t9j h�  h khth@tj
h   ������Q�UR�=�����P�;������} t������������
ǅ���    �����Q�UR�����P�MQ�UR�EP�ݝ����������E������   ��}u�D������Ë�����M�d�    Y_^[�M�3�蠜����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � �����������������������U��Q�E�   ���U�zx t�E�Hx�   ���E���    t�M���   �   ���M�y| t�U�B|�   ���U���    t�E���   �   ���E�    �	�E����E��}�q�M����U�|
��t&�E����M�| t�U����E�L�   ���E����M�| t&�U����E�| t�M����U�D
�   ��뀋U���   �   �   ����]���������������������������������������������������������������������������������U��Q�E���    ��   �M���   (���   �U�zx ��   �E�Hx�9 ��   �U���    t4�E���   �9 u&j�U���   P��������M���   R��������E�x| t.�M�Q|�: u#j�E�H|Q��������U���   P薌����j�M�QxR螇����j�E���   Q芇�����U���    to�E���   �9 uaj�U���   -�   P�W�����j�M���   ��   R�=�����j�E���   ��   Q�#�����j�U���   P�������M���   ��t8�U���   ���    u&�M���   R������j�E���   Q�Ȇ�����E�    �	�U����U��}��  �E����M�|��tR�U����E�| tB�M����U�D
�8 u0j�M����U�D
P�_�����j�M��U����   P�G������M����U�|
 t�E����M�| uF�U����E�| u�M����U�|
 t&h`{hpjj h�   hP}j�Aw������u̋M����U�|
 t:�E����M�| t*�U����E�L�9 uj�U����E�LQ藅���������j�UR脅������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�} �  �E������U�zx t�E�Hx������E���    t�M���   ������M�y| t�U�B|������U���    t�E���   ������E�    �	�E����E��}�m�M����U�|
��t$�E����M�| t�U����E�L������E����M�| t$�U����E�| t�M����U�D
�����넋U���   �   ������E��]������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    襦���E��E��Hp# �t	�U��zl uDj�=u�����E�    �4�P�M���lQ�߶�����E��E������   �j�_��������B����Pl�U�}� u
j 趈�����E�M�d�    Y_^[��]�������������������������������������������������������U��Q�} t�} u3��\�E��M��U�;UtI�E�M��UR�z������}� t�E�P耈�����}� t�M��9 u�}�8�t�U�R胔�����E��]���������������������������������������������U��=�� uj����������   3�]�������������U��Q�E�E��M���  �M��}�wP�U���X��$�D��   k� ���}�1�   �� ���}�!�   �዁�}��   k����}�3���]Ë�����,�<� �����������������������������������������������������U��j�h8d�    P��$���3�P�E�d�    �E�    �E�P�M��{���E�    ���    �}�u)���   ��E��E������M�謋���E��}�c�}�u)���   ��E��E������M��}����E��N�4�}�u.���   �M��g�����Q�U��E������M��G����E���E�E��E������M��-����E��M�d�    Y��]�������������������������������������������������������������������������������U��Q�E�    �	�E����E��}�  }�MM��A ��U�B    �E�@    �Mǁ      �E�    �	�U����U��}�}3��M��Uf�DJ���E�    �	�E����E��}�  }�MM��U���p��A���E�    �	�M����M��}�   }�UU��E���q���  �׋�]���������������������������������������������������������U���   ���3ŉE�������P�M�QR�L���J  ǅ����    ���������������������   s�������������������и   k� Ƅ���� �   k� ������������������������������������tP�����������������������������������B9�����w������   s������Ƅ���� ���j �U�BP������Qh   ������Rjj �J�����j �E�HQh   ������Rh   ������Ph   �M��  Rj �2�����$j �E�HQh   ������Rh   ������Ph   �M��  Rj �������$ǅ����    ���������������������   ��   ��������M������t:�E������H���U������J�E�������������������  �]��������E������t:�U������B�� �M������A�U�������������������  ��U�����Ƃ   �2�����   ǅ����    ���������������������   ��   ������Ar?������Zw6�M������Q���E������P�������� �U�������  �X������ar?������zw6�E������H�� �U������J�������� �M�������  ��U�����Ƃ   �<����M�3�������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hКh�Ld�    P���SVW���1E�3�P�E�d�    �E�    �u����E��E��Hp# �t�U��zl ��   j�	l�����E�    �E��Hh�M�U�;|�tK�}� t$�E�����Iu�}�X�tj�U�R�py�����E��|��Hh�|��U�E�   ���E������   �j��������	�U��Bh�E�}� u
j �=�����E�M�d�    Y_^[��]������������������������������������������������������������������������������U����E�    �E�P�M���s���M������H�y t �M������P�B�E��M������E����E�    �M��ԃ���E���M��ǃ����]���������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�����腛���E�耧���E܋Hh�M��UR�*������E�E��M;H�  h[  h�}jh   �e�����E��}� ��  �Uܹ�   �rh�}��E��     �M�Q�UR�j�����E؃}� ��  �E܋Hh�����Ju�E܁xhX�tj�M܋QhR�5w�����E܋M��Hh�U܋Bh�   ���U܋Bp���1  � ����"  j�Ii�����E�    �U��B����M��Q����E���  ����E�    �	�U���U�}�}�E�M�U�f�LJf�E�����E�    �	�U���U�}�  }�E�E�M�P��P����E�    �	�E���E�}�   }�M�M�U䊁  ��X��׋|������Ju�=|�X�tj�|�P�v�����M��|��U�   ���E������   �j苠������(�}��u"�}�X�tj�M�Q�u�����y����    ��E�    �E؋M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���,���3ŉE�V�EP�&������E�} u�MQ�a�����3��0  �E�    �	�Uԃ��Uԃ}��t  kE�0����;M�\  �E�    �	�U���U�}�  s�EE��@ ���E�    �	�M����M��}���   kU�0�E�����M��	�U܃��Uܸ   k� �U��
��ts�   �� �U��
��t`�   k� �E���M��	�U���U�   �� �M��9U�w*�}�   s!�E���x��UU��B��MM�A��q����F����U�E�B�M�A   �U�BP��������M��  �E�    �	�U����U��}�skE�0�M��U�u�f��p��f�DJ�ՋMQ�������3��  �y����} t!�}��  t�}��  t�UR� ��u����q  �E�P�MQ�L���?  �E�    �	�U���U�}�  s�EE��@ ��M�U�Q�Eǀ      �}���   �M�M��	�U؃��U؋E����tE�U��B��t:�M���U��	�E���E�M��Q9U�w�EE��H���UU�J����E�   �	�E���E�}��   s�MM��Q���EE�P�֋M�QR�|������M��  �U�B   �
�E�@    �E�    �	�M����M��}�s3ҋE��Mf�TA��UR�Z�����3���=�� t�EP�1�����3�����^�M�3�虁����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��}�|	�}�   ~#h�}hpjj j8h0~j�a������u̋MQ�URj �s]����]������������������������U����EP�M��<k���}�|	�}�   ~#h�}hpjj jDh0~j�Ea������u̃}�|5�}�   ,�M��K�������   �M�H#U�U��M��%{���E��9�/�M������ �   k�����   �#M�M��M���z���E���M���z����]�������������������������������������������������������U��=4� u�E����A#E��j �UR�EP�t����]�����������������������������U���0�EP�M���i���}�|6�}�   -�M��=�������   �E�B#M�M�M��z���E���   �M�����P�U�����   R��������tN�E��%�   �   k� �D��   �� �M�L��   ��U�}�s��m����E��D� �E�   �2�   k� �E�D��E�   �}�s��9����M��D� �E�   j�M��l�����BP�M�Q�U�R�E�Pj�M��P���P��������u�E�    �M��+y���E���M�#M�M��M��y���E���]�������������������������������������������������������������������������������������������������U��QV�E�    �} u�4�EPj ���Q��E��}� u��P�O�������賤���0^��]��������������������U���V�E�E��} u�MQ膂������   �} u�UR視����3��   �E�    �}�w)�} u�E   �EP�MQj ���R��E���EP�5����������    3��e�}� u	�=�� u%�}� t���P�z��������ޣ���0�E��1�MQ��������u��P�M�������豣���03���J���^��]�������������������������������������������������������������������������U���V�} t	�E�   ��E�    �E��E�}� u#h�~hpjj jLh�~j�\������u̃}� u-�����    j jLh�~h h�~�P�����3��   �}�v�Ϣ���    3��~�} u�E   �URj ���P��E��MQ�URj���P��E��}� u:�}� @  w�M;M�w�u   ��t�U�U����P���������L����0�E�^��]��������������������������������������������������������������������������U����E�����j j�E�Pj ���Q���t�}�u	�E�   ��E�    �E���]����������������������������U����E�E��M�Q�UR�EP�MQ�UR�EP�MQ��Z�����E��E�    �E���]��������������������������������U��E P�MQ�UR�EP�MQ�UR�EP萔����]������������������������U��j�h@�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t�}t	�E�    ��E�   �E܉E؃}� u#h��hpjj jth�j�Z������u̃}� u.�l����    j jth�hTh��躘��������  �} t	�E�   ��E�    �UԉUЃ}� u#h��hpjj juh�j�Y������u̃}� u.�����    j juh�hTh���A���������  j�TZ�����E�    �T��M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���M̋U�ẺB�M̉M��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H�T�j�U�R�Wg�����<3�u&h��hpjj h�   h�j�X������u��E������ߞ���    ��   �}� tu�U�B���EȋM�UȉQ�EȉE��M�;T�tM�U�z t�E�H�U���M��E�H�J�U��    �E�T��H�T��E��M�T��h�   h<�jj��S�����E�}� u�E������.����    �L�U��    �E�T��H�=T� t�T��E��M��A   �E�   �U�E�B�M�T��E������   �j诐����ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��X!  �R������3ŉE�ǅ����    ǅ����    ǅ����    �} u
�   �N  ������P�MQj�,��u
ǅ����    �   i�  ������������  s������������Ƅ���� h  ������R������P���u8j h_  h�h�h�h4�h  ������Q�.�����P�b`����������������������P�������@vl������Q�}�����������D�������j hh  h�h�hX�j�x�Q������������+й  +�Q������R�a����P��_�����} t*�EP�������@v�MQ��~�����U�DÉ������+���������������     �}uǅ����h��
ǅ����p��   k� �M���t�E�������
ǅ�����a�   k� �E���t�}uǅ����|��
ǅ����p��   k� �M���tǅ�������
ǅ����p��} t�E�������
ǅ�����a�} tǅ�������
ǅ����p��} t�M�������
ǅ�����a�} tǅ�������
ǅ����p������� t�������������'�} t�E�������
ǅ�����a������������������ tǅ����t��
ǅ����p��} tǅ�������
ǅ����p�������R������P������Q������R������P������Q������R������P������Q������R������P������Q�U��@PhP�h�  h   ������Q�u����D������������ }*j h  h�h�h��j"j�����R��O���� �ژ��������������� }8j h�  h�h�h��h��h   ������R�t�����P�]����h  h��������P�q����������������uj�`����j��S��������u�   �3��M�3��p����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��|�]�������U��� ]������U���D]������U��j�h`�h�Ld�    P���SVW���1E�3�P�E�d�    �E�E�}� ��  �M�y$ tj�U�B$P�^�����M�y, tj�U�B,P�^�����M�y4 tj�U�B4P�^�����M�y< tj�U�B<P�q^�����M�y@ tj�U�B@P�W^�����M�yD tj�U�BDP�=^�����M�yH tj�U�BHP�#^�����M�y\��tj�U�B\P�^����j�PP�����E�    �M�Qh�U܃}� t$�E܃����Iu�}�X�tj�U�R��]�����E������   �j�W������j��O�����E�   �E�Hl�M��}� t4�U�R��c�����E�;4�t�}�8�t�M��9 u�U�R��o�����E������   �j�������j�E�P�.]�����M�d�    Y_^[��]� ���������������������������������������������������������������������������������������������������������������������������������U��=|��t1�} u�|�P��f�����Ej �|�Q�W�����UR�O���]������������������U��Q�����E��}� u
j�Ob�����E���]��������������U������E��|�P�Vf�����E��}� uwj h  h,�jh�  j�u�����E��}� tQ�M�Q�|�R�W������t%j �E�P�dc�����D�M���U��B�����j�E�P�[�����E�    �M�Q�X�E���]���������������������������������������������������U��j�h��h�Ld�    P��SVW���1E�3�P�E�d�    �E�@\���M�A    �U�B   �E�@p   �   k� �C   �Mf���   �   k� �C   �Uf���  �E�@hX��Mǁ�      j��L�����E�    �U�Bh�   ���E������   �j�������j�L�����E�   �U�E�Bl�M�yl u�U�4��Bl�M�QlR�_�����E������   �j蹄����ËM�d�    Y_^[��]���������������������������������������������������������������������������������U��Q�Ԛ��輊����u�8~��3��   h<\��[�����|��=|��u	�~��3��ijrh,�jh�  j�'c�����E��}� t�E�P�|�Q�T������u	��}��3��(j �U�R��`�����D�M���U��B�����   ��]��������������������������������������������������U��=|��t�|�P�w�����|�������h��]����������������������U����P�]����������������U��} t#h`�hpjj jWhx�j�I������u�j �h����]�������������������������U��Qj�_J�������P��E��MQ����j萂�����E���]��������������������U��Q���P��E��}� t�MQ�U�����u3���   ��]�����������������������������U��E���]����U��Q�E�����j j ���P�0��u�E������E���]��������������������U���q��]�������U��Q�=�� u�P���j�Ar����h�   �r�����} t�E�E���E�   �M�Qj ���R�$��]����������������������������U��Q�E�    �}�wC�EP�f�����E��}� t�*�=�� u�3����    ��MQ�:�������u����UR�$����������    3���}� u�����    �E���]������������������������������������������U��=�� u#hȅhpjj jXh��j�*G������u̡��]���������������������������U���(����=�� u3���   ]���������������U�����    ]������������������U���SQ�E���E��EU�u�M�m��cR��VW��_^��]�MU���   u�   Q�AR��]Y[�� ��������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �e���P��E�}� t#�E�    �U��E�������   Ëe��E������G���M�d�    Y_^[��]�����������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �e��w���@x�E�}� t#�E�    �U��E�������   Ëe��E������c���M�d�    Y_^[��]�����������������������������������U��Q�8w���@|�E��}� t�U��F����]����������������U��hv'����]������������U��j�h �h�Ld�    P���SVW���1E�3�P�E�d�    �E�x �Q  h (  hI^hJj �M��	Qj ��w�����E��}� u3��%  �U�R�^n�����E�E�EԋM���M�}� v�U�U���� u�M�M�� ��j��D�����E�    �U�z ��   j�Qh�����E܃}� ��   �E��P�5h�����E؋M�U؉Q�}� t[j h�   hx�h؆h��E�P�M��Q�U�BP� �����P�TN�����M܋U�B��M܋U�B�A�M�U܉Q��E�P��{�����M�Q��{�����E������   �j�y|����ËU�B�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������U��j�h@�h�Ld�    P���SVW���1E�3�P�E�d�    �E�x �f  j�VC�����E�    �M�y �/  h (  j �U��	Rj �'������E��}� u"�E�    j��E�Ph���F������E��  �M�Q�l�����E�U�UЋE���E�}� v�M�M���� u�E�E��  ��j�0f�����E܃}� ��   �E�    �M��Q�f�����E؃}� taj h  hx�hȇh��U�R�E��P�M�Q������P�8L�����U�E؉B�M܋U�B��M܋U�B�A�M�U܉Q��E�P��y�����M�Q��y�����E������   �j�Tz����ËU�B�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������U��j�h �h�Ld�    P���SVW���1E�3�P�E�d�    j�3A�����E�    �E�x ��   ����M��E�����U��U�}� t[�E�M�;Qu�E��M�Q�P�E�P�x�����4�M�M��U�z u#hD�hpjj j9hx�j�?������u�뙋M�QR�Fx�����E�@    �E������   �j��x����ËM�d�    Y_^[��]����������������������������������������������������������������������U��j�h`�h�Ld�    P���SVW���1E�3�P�E�d�    j��?�����E�    �E�x ��   ����M��E�����U��U�}� t^�E�M�;Qu�E��M�Q�P�E�P�;w�����7�M�M��U�z u&hD�hpjj h�   hx�j�a>������u�떋M�QR��v�����E�@    �E������   �j�{w����ËM�d�    Y_^[��]�����������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    j�>�����E�    �E�H�M��E�    ��U��U�}� t%�E�H�M��U�P��u�����M�Q��u�������E������   �j�zv����ËM�d�    Y_^[��]��������������������������������������������������U���E��u	� (  f�M�URhI^hJ�EP�MQ�UR�<p����]������������������������U��EP�MQ资����]������������U��j �EP�MQ�UR�EP�MQ�UR�XZ����]����������U��Q�E�    �}et�}Eu%�E P�MQ�UR�EP�MQ�UR�7�����E��{�}fu!�E P�MQ�UR�EP�MQ�������E��T�}at�}Au%�U R�EP�MQ�UR�EP�MQ�x6�����E��#�U R�EP�MQ�UR�EP�MQ蝂�����E��E���]���������������������������������������������������U��j �EP�MQ�UR�EP�MQ��5����]��������������U���   �E�E��E��  �E�    �E�    �E�    �0   f�M��E�    �E�    3�f�U��E�    �E�    �E�    �E�    �EP��X����{D���} }�E    �} t	�E�   ��E�    �M��M��}� u&h��hpjj h�  h��j�a:������u̃}� uI趀���    j h�  h��hЊh���y����ǅh���   ��X����1T����h����L  �} v	�E�   ��E�    �E��E��}� u&h�hpjj h�  h��j��9������u̃}� uC�����    j h�  h��hЊh��jx�����E�   ��X����S���E��  �   k� �M� �U��9Uv	�E�   ��E�    �E��E��}� u&h�hpjj h�  h��j�%9������u̃}� uI�z��� "   j h�  h��hЊh���w����ǅt���"   ��X�����R����t����  �U܋�R�4�rR��%�  �� �E��U��}��  �  �}� �  �}�u�E�E��	�M���M�j �UR�E�P�M��Q�UR��@�����Eȃ}� t(�   k� �U�
 �EȉE���X����YR���E��w  �   ��U�
��-u�M�-�U���U�E� 0�M���M�} t�E�X��E�x�U�E��M���Mje�UR��a�����E��}� t'�} t�E�P��E�p�E��M��U����U��E��  �MȉM���X����Q���E���  �U܋�R�?�0Q������ �E��U��E�E�t�M�-�U���U�E� 0�M���M�} t�E�X��E�x�U�E��M���M�} t�E�A��E�a�U��:�UċM܋�Q�4�P��%�  �� �E��U��U�U�u[�E� 0�M���M�U܋�J���� ��x�����|�����x����|���u�E�    �E�    ��Ẽ��MЃ� �ẺM���U�1�E���E�M�M��U���U�} u�E��  ���X����~�������   ��M����E܋�P���� ��l�����p�����p��� w��l��� �p  �E�   �E�    �M�EԋU��Ƃ���EԉU��E����   �} ~}�M܋�Q���� #E�#U��M��yO��f�E��U���0f�U��E���9~�M�M�f�M��U�E���M���M�EԋUر�8O���EԉU��U��f�U�E���E�q����M����   �U܋�R���� #E�#U��M���N��f�E��E�����   �M�M��U����U��E����ft�U����Fu�M��0�U����U��ًE�;E�t/�M����9u�E���UčD�M����U�����M����U����U��E�����U��
�	�E���E�} ~�M�0�U���U���E����u�U��U�} t�E�P��E�p�E�M��U���U�M܋�Q�4��M��%�  �� +E�UЉE��U�}� |�}� r�U�+�E���E�"�M�-�U���U�E��؋M�� �ىE��M�U�U��E�� 0�}� |M	�}��  rBj h�  �M�Q�U�R�l�������0�M��U���Uj h�  �E�P�M�Q�����E��U�U;U�u�}� |D�}�dr<j jd�E�P�M�Q�����Ѓ�0�E��M���Mj jd�U�R�E�P�ʀ���E��U�M;M�u�}� |D�}�
r<j j
�U�R�E�P�ŀ���ȃ�0�U�
�E���Ej j
�M�Q�U�R�x����E��U��E���0�M��U���U�E�  �E�    ��X�����L���E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�EP�MQ�+����]��������������U���\�E�    �E P�M��%:���} t	�E�   ��E�    �M��M�}� u&h��hpjj h�   h��j�0������u̃}� u@�mv���    j h�   h��h�h���n�����E�   �M���I���E��\  �} v	�E�   ��E�    �E�E�}� u&h�hpjj h�   h��j�/������u̃}� u@��u���    j h�   h��h�h��*n�����E�   �M��`I���E���  �} ~�U�U���E�    �E���	9Ev	�E�   ��E�    �M܉M؃}� u&hH�hpjj h  h��j��.������u̃}� u@�7u��� "   j h  h��h�hH��m�����E�"   �M��H���E��&  �E��tG�M�9-u	�E�   ��E�    �UUԉU��} ~	�E�   ��E�    �E�P�M�Q�w  ���U�U��E�8-u�M��-�U����U��} ~-�E��M��Q��E����E��M��+{������   ��M����E��t	�E�    ��E�   �M�MM̉M��}�u�U�U���E�+E�M+ȉM�j h%  h��h�h؉h���U�R�E�P�+u����P�_8�����M����M�} t�U��E�E����E��M�Q���0��   �M�Q���U�y�E��؉E��M��-�U����U��}�d|)�E���d   ���ЋE��ʋU��
�E���d   ���U��U����U��}�
|)�E���
   ���ЋE��ʋU��
�E���
   ���U��U����U��E��M��ЋE��� ���t �U����0uj�M��Q�U�R�5�����E�    �M��F���E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���\���3ŉE��E�E��M��M��E�    j�U�R�E�P�M��QR�P�W>�����} t	�E�   ��E�    �M��M��}� u&h��hpjj hn  h��j��*������u̃}� u3�7q���    j hn  h��h��h���i�����   �]  �} v	�E�   ��E�    �E��Ẽ}� u&h�hpjj ho  h��j�a*������u̃}� u3�p���    j ho  h��h��h��i�����   ��   �}�u�U�U��:�E܃8-u	�E�   ��E�    �} ~	�E�   ��E�    �M+M�+MĉMԋU܃:-u	�E�   ��E�    �} ~	�E�   ��E�    �E�P�M��Q�U�R�EE�E�P�F�����E��}� t�   k� �E� �E��(�MQj �U�R�EP�MQ�UR�EP��������E��E��M�3��H����]������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�EP�n����]������������������U���@�E�H���M��UR�M�� 2���} t	�E�   ��E�    �E�E��}� u&h��hpjj h�  h��j�(������u̃}� u@�hn���    j h�  h��hL�h���f�����E�   �M���A���E���  �} v	�E�   ��E�    �U�U�}� u&h�hpjj h�  h��j�'������u̃}� u@��m���    j h�  h��hL�h��%f�����E�   �M��[A���E��R  �M��tG�U�:-u	�E�   ��E�    �EE�E��M�;Mu�U�U��U��E�� 0�M����M��U�� �E�E��M�9-u�U��-�E����E��M�y j�U�R��
  ���E�� 0�M����M���U�E�B�E��} ��   j�M�Q�
  ���M��s������   ��U����M����M��U�z }]�E��t�M�Q�ډU�&�E�H��9M}�U�U���E�H�ىM܋U܉U�EP�M�Q�;
  ���URj0�E�P�	M�����E�    �M��@���EЋ�]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���T���3ŉE��E�E��M��M��E�    j�U�R�E�P�M��QR�P�'8�����} t	�E�   ��E�    �M̉Mă}� u&h��hpjj h�  h��j�$������u̃}� u3�k���    j h�  h��hd�h���Rc�����   �*  �} v	�E�   ��E�    �E��E؃}� u&h�hpjj h�  h��j�1$������u̃}� u3�j���    j h�  h��hd�h���b�����   �   �}�u�U�U��!�E܃8-u	�E�   ��E�    �M+MȉMԋU܃:-u	�E�   ��E�    �E�P�M܋UQR�E�P�MM�Q�@�����E��}� t�   k� �M� �E��$�URj �E�P�MQ�UR�EP��������E��E��M�3��	B����]�����������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�EP�MQ�i����]��������������U���d���3ŉE��E�    �E�E��E� �M��M�j�U�R�E�P�M��QR�P�s5�����} t	�E�   ��E�    �MĉM��}� u&h��hpjj h-  h��j��!������u̃}� u3�Sh���    j h-  h��h|�h���`�����   �  �} v	�E�   ��E�    �ẺE��}� u&h�hpjj h.  h��j�}!������u̃}� u3��g���    j h.  h��h|�h��`�����   �9  �U܋B���EԋM܃9-u	�E�   ��E�    �UU��U؃}�u�E�E��!�M܃9-u	�E�   ��E�    �U+U��UȋE�P�MQ�U�R�E�P��=�����EЃ}� t�   k� �E� �E��   �M܋Q��9U�}�E���E� �E�E�M܋Q���Uԃ}��|�E�;E|&�MQj�U�R�EP�MQ�UR�EP��������I�G�M��t!�U���E��M؃��M؃}� t��U��B� �EPj�M�Q�UR�EP�MQ�������M�3���>����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�aF����]��������������U���V�EP�M���(���M���t*�E�0�M��+l������   ��;�t�U���U�̋E��M��U���U�}� ��   �E���t!�U���et�M���Et�E���E�ՋM�M��U���U�E���0u�U���U��E�0�M��k������   ��;�u	�U���U�E���E�M�U����M��U�E����E��}� t�ӍM��=8��^��]����������������������������������������������������������������������������U��j �EP�MQ�UR��b����]����������������������U����} t$�EP�MQ�U�R�|G�����E�M��U��P��EP�MQ�U�R��Q�����E�M����]���������������������������������U��j �EP��1����]��������������U����EP�M���&���M�R�VY������et�E���E�M�R�j������u�E�Q�&Y������xu	�U���U�E��M��M���i������   ��U���M���M�U��E��M�U���E��E��M��U��E���E�}� uҍM��n6����]��������������������������������������������������������������U��Q�E�������Az	�E�   ��E�    �E���]������������������������U��} t#�EP��E������P�MQ�UUR�D$����]�������������������U��j jh��h�h8�h   h   j �I,����P�<&����]����������������������������U��Q�E�    �	�E����E��}�
s�M���0�R��M���0��ԋ�]��������������������U����Te���E��}� u3���  �E��H\Q�UR�  ���E��}� u	�E�    �	�E��H�M�}� u3��  �}�u�U��B    �   �  �}�u����t  �E��H`�M�U��E�B`�M��y�2  �H��U��	�E����E��H�L�9M�}kU��E��H\�D    �ҋU��Bd�E�M��9�  �u�U��Bd�   �   �E��8�  �u�M��Ad�   �   �U��:�  �u�E��@d�   �   �M��9�  �u�U��Bd�   �q�E��8�  �u�M��Ad�   �Z�U��:�  �u�E��@d�   �C�M��9�  �u�U��Bd�   �,�E��8� �u�M��Ad�   ��U��:� �u
�E��@d�   �M��QdRj�U���E��M�Hd��U��B    �E��HQ�U���U��E�B`�����]�������������������������������������������������������������������������������������������������������������������������������������������U��}csm�u�EP�MQ�y-������3�]�������������U��Q�E�E��M��;Ut�E����E�k@�M9M�s��k@�U9U�s
�E��;Mt3���E���]�������������������������������U��E�(�]����U����E�    �=�� u�7���   i�  �M��}�  s��aV���U�Ƃ�� h  h��j �h����7�����=H� t�H����t�H��U���E����E�E�M�Q�U�Rj j �E�P��   ���}����?s�}��r����w�M��U���;E�s����dh�   hp�j�M��U���P�������E�}� u����8�M�Q�U�R�E��M��R�E�P�M�Q�w   ���U������E���3���]�������������������������������������������������������������������������������������������U��� �E�     �M�   �U�U��} t�E�M��U���U�E�    �E����"u/�}� u	�E�   ��E�    �U�U��E���M��U����U��w�E����U�
�} t�E�M����E���E�M���U��E����E��M�Q�W#������t/�U����M��} t�U�E���
�U���U�E����E��M���t �}� �=����U��� t�E���	�'����M���u�U����U���} t�E�@� �E�    �M����t!�E���� t�U����	u�M����M��ߋU����u��  �} t�M�U��E���E�M����E��E�   �E�    �M����\u�E����E��M���M���U����"u`�E�3ҹ   ���uH�}� t�   �� �E����"u�U����U��#�E�    �}� u	�E�   ��E�    �E�E��M���M�U�U��E���E�}� t$�} t�M�\�U���U�E����U�
�ǋE����t�}� u�U���� t�M����	u�   �}� ��   �} tQ�E��Q�\!������t)�U�E���
�U���U�E����E��M����E��M�U����M���M�)�U��P�!������t�M����M��U����M��U����M��U����U��_����} t�E�  �M���M�U����M�������} t�U�    �E���E�M����E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����=�� u�1���E�    ����E��}� u����e  �M����t,�E����=t	�U���U�E�P�;�����M��T�U���juh��jj�E��P��)�����E��M�� ��= � u�����   ����U��	�E�E��E��M������   �E�P�;�������E��M����=��   j~h��jj�E�P�I)�����M���U��: uj� �P�T����� �    ����rj h�   h؍h@�hX��M�Q�U�R�E��Q�X����P�F�����U����U��B���j���P���������    �M��    ���   3���]�������������������������������������������������������������������������������������������������������U����E�    �E�    �=��N�@�t���%  ��t����щ���   �U�R�4�E�E��M�3M��M��D3E��E��03E��E��U�R�,�E�3E�E��M�3M��M��U��E�3ЉU��}�N�@�u	�E�O�@���M���  ��u�U���G  ��U��U��E�����M��щ����]��������������������������������������������������������������������U����E�    �8�E��}� u3���   �E��E��M����t�E����E��M����u	�E����E��؋M�+M������M�j j j j �U�R�E�Pj j ��E��}� tjJh��j�M�Q�
�����E�}� u�U�R�<3��Dj j �E�P�M�Q�U�R�E�Pj j ���uj�M�Q�k�����E�    �U�R�<�E��]���������������������������������������������������������������������������V�E��=�Gs����t�Ѓ����Gr�^������������V��H��=Ks����t�Ѓ���Kr�^������������U��EPj �MQ�UR�EP�IO����]������������������U���@�E�    3��EĉEȉẺEЉEԉE؉E܍M��M��} t	�E�   ��E�    �U��U�}� u#h��hpjj jphȎj�j������u̃}� u.�R���    j jphȎh,�h���K��������.  �} t�} u	�E�    ��E�   �M��M�}� u#hP�hpjj jshȎj��������u̃}� u.�@R���    j jshȎh,�hP��J��������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R�}C�����E�} u�E��P�E��H���M�U��E�B�}� |!�M��� 3�%�   �E��M�����E����M�Qj �ZJ�����E��E��]���������������������������������������������������������������������������������������������������������������������������̀zuf��\���������?�f�?f��^���٭^�������剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�������剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp���������۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-����p��� ƅp���
��
�t�������������������������������������������������������������������������������������������������������������������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�:�����E�f�}t�m���������������������������������������������������ËT$��   ��f�T$�l$é   t�   �����   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   ����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t���Z��9��Z��,$Z���������������������   s�����������������������   v��������������������������������������������������������������������������������������������������������U��Q�E�   �} u�E�    �E���]������������������U��Q�E�   �} u�E�    �E���]������������������U��Q�E�   �} u�E�    �E���]������������������U��3�]����������U��j�h@�h�Ld�    P��SVW���1E�3�P�E�d�    �=4�8�tAj�������E�    h8�h4��G�����4��E������   �j�>����ËM�d�    Y_^[��]��������������������������������������������������U��@�]�������U��0�]�������U����} u3��   jU�EP�A�����E��}�Ur3��ihw  hĒj�M��T	R�' �����E��}� u3��@j hz  h0�h̤h ��E���P�MQ�U���R�E�P�����P������E���]������������������������������������������������������U��EP�MQ�9����]������������U��EP�����]����������������U���m��]�������U��j hc  h0�h �h@��EP�MQ�UR�VJ����P�������   k� �U��
�   ��t!�M���   QhĤj�UR�EP�_(�����   k� �E��   ��t!�U��   RhȤj�EP�MQ�'(����]���������������������������������������������������������U���h�  j �EP�Z)�����M���u3���  �   k� �U�
��.up�   �� �U�
��t]j h9  h0�h�h0�j�   �� MQj�U��   R�����P������   k�3ҋEf��   3��j  �E�    �	�M���M�h4��UR�I�����E��}� u����6  �E��Mf�Af�U��}� uI�}�@sC�E���.t:j hG  h0�h�h@��M�Q�URj@�EP������P������   �}�uL�}�@sF�M���_t=j hJ  h0�h�h8��U�R�EPj@�M���   Q�����P������^�}�uS�}�sM�U���t	�E���,u<j hM  h0�h�h(��M�Q�URj�E   P�@����P�W���������)�M���,u��U���u��E��M�TA�U����3���]�����������������������������������������������������������������������������������������������������������������������������������������������������U�����1���E��E��Hp��u	�E�   ��E�   �U�U�E�E��M����M��}�wC�U��$��&�E��Hp���U��Jp�   �E��Hp����U��Jp�   �   � ������z3�t	�E�   ��E�    �M��M�}� u&h��hpjj h�   h0�j���������u̃}� u.�AE���    j h�   h0�h��h���=���������E��]�k&f&>&R&������������������������������������������������������������������������U��VW�} t0�} t*�E;Et"�.   �u�}�M�    �UR�'����_^]������������������U���  ���3ŉE��} |�}�} u3��7h�   ������Pj��MQj j ���u3��������R�EP�-2�����M�3��c����]�����������������������������������U���  ���3ŉE��/���   ��(�����(������� �����(����������ǅ����   ��(�����"  ��$���ǅ����   ǅ,���    ǅ���    �} u3��T  j h�  h0�hT�hx�jU��(���P  P�MQ�UR�s����P������E���Cu^�   �� �E���uKj h�  h0�hT�h�hp��UR�EP�C����P�8�����} t	�M�    �E�  �UR��%������,�����,����   s6�EP��$���Q�&�������  �UR�����P�e&�������  ǅ����p�ǅ ���    ǅ���    ǅ���   �   k�����3�������t
ǅ���    �MQ��0���R�f4������uQ����� t%��0���P�� ���Q��0���R�^&����������#��0���P�� ���Q��0���R��$�������������� tq��0���P�����Q��$���R�J�����} tIj h�  h0�hT�hx���P���P�$������P��P���Q�UR�EP�����P������m  �MQ�uD�������  j�����Rh  �EP��������t	����� u������������� ����
j h�  h0�hT�hp���,�����P�MQ�����R��$���P������P�����j h�  h0�hT�h���,�����Q�UR�EP�MQ�����P������j h�  h0�hT�h����,�����R�EPjU��(�����P  Q�l����P������Qj h  h0�hT�hp��UR�1#������P�EPjU��(�����P  Q� ����P�7����3��   �U���tQ��,����   sEj h  h0�hT�h ���,�����Q�UR�����P�����Q������P�������3ҋ����f��} tj�� ���Q�UR�����j h  h0�hT�h����$���P�MQ�UR��?����P�y������$����M�3��W����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hМh�Ld�    P��SVW���1E�3�P�E�d�    �} ��   j��������E�    �E�x t-�M�Q�����Hu�M�yX�tj�U�BP�h�����E������   �j��/����ËM�9 tcj�������E�   �U�P������M�9 t#�U��8 u�M�98�t�U�P������E������   �j�/�����j�MQ�������M�d�    Y_^[��]����������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    ��'���E�h�  hĒjjj�������E�}� u��;���    3��   �P0���3���E�M��Ql��E�M��Qh�Pj�0������E�    �E�Q�0	�����E������   �j�\.�����j��������E�   �U�B�   ���E������   �j�#.����ËE�M�d�    Y_^[��]������������������������������������������������������������������������U����E�    �} |�}�} u3��  hL  hĒjjj������E��}� u�:���    3��  hQ  hĒjjh�   �}�����E��E��M���}� u j�U�R������A:���    3��=  hW  hĒjjh   �1�����E�E��M�H�}� u0j�U��P�7����j�M�Q�)������9���    3���   h8��U��P�������MQ�UR�E��Q�x	  ����uDj�U��BP�������M��R�L�����E��Q�d����j�U�R������E�    �l�E��HQ�U���HQ�<�������tDj�U��BP�y�����M��R�������E��Q�����j�U�R�O�����E�    ��E��H�   �E���]���������������������������������������������������������������������������������������������������������������������������U����E�E��E�    �	�M����M��U�;U}A�E����E�j h&  h0�h �h8��M��Q�R�EP�MQ��9����P��������E�    ��]�������������������������������U��j�h �h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} |�}	�E�   ��E�    �E؉Eԃ}� u&h��hpjj h  h0�j���������u̃}� u0�R7���    j h  h0�h`�h���/����3��  ��"���E��+���U��Bp���M��Ap�E�    h  hĒjjh�   �	�����E�}� �  j�f������E�   �U��BlP�M�Q�������E�    �   �j�)����Ã}� ��   �UR�EP�M�Q�K  ���E܃}� ��   �} th���UR�c������t
�4�   j��������E�   �E�P�M���lQ�}2�����U�R�������E��Hp��u$� ���u�E��HlQh4��G2�����g  �E�    �   �j��(�������U�R������E�P������E������   ��M��Qp���E��PpËE܋M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�   �E�    �E�    �E�    �E�    �E�  hd  hĒj�E�P�I������E�}� u3��X  �M���M��U�����U�3��M�f��U��   �E�   �	�E����E��M����U�D
Ph�kM���8�Rj�E�P�M�Q�N�����}�}kj hp  h0�h�h�h���U�R�E�P�5����P�f������M������U�D
P�M����U�D
P��������t�E�    �{  �}� �/  �   k� �E�| tZ�   k� �E�L�����JuA3�u#j hpjj hy  h0�j���������u�j�   k� �M�TR�������   k� �U�|
 tZ�   k� �U�D
�����IuA3�u#j hpjj h~  h0�j��������u�j�   k� �E�LQ�������   k� �M�D    �   k� �M�D    �   k� �M�U�T�   k� �U�E��D
�E��L  �B  j�M�Q�������   k� �M�| tZ�   k� �M�T�����HuA3�u#j hpjj h�  h0�j���������u�j�   k� �U�D
P�F������   k� �E�| tZ�   k� �E�L�����JuA3�u#j hpjj h�  h0�j�T�������u�j�   k� �M�TR��������   k� �U�D
    �   k� �U�D
    �   k� �U�D
    �   k� �U�D
    �   ���M�D��������]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����  ���3ŉE��} tF�} t�EP�MQ�UR�0  ����,�����E���M�T��,�����,�����0�����  ǅ ���   ǅ4���    �} ��  �   k� �E���L�a  �   �� �E���C�I  �   ��E���_�2  �U��<���h|���<���P��$������@�����@��� t$��@���+�<�������8���t��@������;u3��  ǅD���   ���D�������D�����D���J��8���R��<���Pk�D�����8�R��0������u k�D�����8�Q�����9�8���u�랋�@�������@���h����@���P�*0������8�����8��� u��@������;t3��f  ��D�����   j h�  h0�h��h����8���P��@���Qh�   ������R�z�����P��������8�������$�����$���  s��k&��3ɋ�$���f������������P��D���Q�UR��  ����t��4�������4�����8�����@����J��<�����<������t��<�������<�����<������������4��� t�EP������������
ǅ���    �������0����&  j jU��H���Rh�   ������P�MQ�d(������0�����0��� ��   ǅD���    ���D�������D�����D���|��D��� tn��D������M�TR������P��������t;������Q��D���R�EP��  ����t��4�������4����
ǅ ���    ���4�������4����l����� ��� t�EP�r�������0����3��4��� t�MQ�U�������(����
ǅ(���    ��(�����0�����EP�)�������0�����0����M�3��]����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����  ���3ŉE�Vǅ<���    ǅ4���    ǅ$���    �z�������������  ��D���ǅ(���   �� ���QjU��H���Rh�   ������P�MQ�%������u3��<  �U���E�LQ������R�7������u�E���M�D�	  ������R�T��������$���h�  hĒj��$����L Q��������<�����<��� u3��  ��<�������4����E���M�T������E�M����   ������E�H�����j h�  h0�hT�h��������R��$���P��4���Q�4*����P��������U���E��4����L�   k� ��������Cu'�   �� ��������u�M�UǄ��       ���H���P�3
�����M�U����   �}�:  �E�� ����H��(�����D����L���T����,�����0���ǅ@���    ���@�������@�����@���;�(�����   �U��@�����D����R;�uT��@��� tG��@�����D������D��   k� ��D�����D��@�����D�����,����Ћ�0����L��]�V��@�����D����ЋT�������������@�����D�����,�������0����T��������,����������0���������@���;�(�����   j�E�HQ������Rjh �jj ����������   ǅ8���    ���8�������8�����8���s$��8�����M�������  ��8���f��E������h�   �`�Q������R���������u�   k� ��D����D
   ��   k� ��D����D
    ��   k� ��D����D
    �   k� ��D����E�@�
�   k� �E��D����T�Pp�&�}u�E�� ����H��}u�U�� ����B�MQkU��@��Ѓ���tb�M���U������D
j�M�U����   P�z������M�U���������   j��<���Q�V������U������B3���   ���������   �M���U�D
�����I��   3�u#j hpjj hH  h0�j�Q�������u�j�M���U�D
P�������j�M���U�D
P�������j�M�U����   P�������M���U�D
    �E�MǄ��       ��<��� t��<����   �E���M��<����T�E���M�D^�M�3��k�����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��4����   � ��4����   ���4��Qt���]���������������������������U����E�    �} u�E��Q�U�}  t	�E�	   ��E�   j j �EP�MQ�U�R�EP��E��}� u3���   3�uS�}� ~M�}����wD�U���R���������t#h��  �E��L Q�u����P������E���E�    �U��U���E�    �E�E��}� u3��a�M���Qj �U�R������E�P�M�Q�UR�EPj�MQ��E�}� t�UR�E�P�M�Q�UR��E�E�P�x������E��]��������������������������������������������������������������������������������U����EP�M������M Q�UR�EP�MQ�UR�EP�M��D(��P�H������E��M��'����E���]��������������������U��EP�MQ�UR�EP�w	����]��������������������U���T�E�    �} t�} u3��`  �} t�} v3��Mf��} t	�E�   ��E�    �U��U�}� u#h|�hpjj jEh��j�P�������u̃}� u.� ���    j jEh��h�h|������������  �MQ�M�������} �  �M��'����   �����    uj�M�;MsG�UU�f��Mf��UU����u�M��M�M�������E��g  �U����U��E���E뱋M��M�M������E��=  �  �UR�EPj��MQj	�M��&����BP��E��}� t�M����M��M��W����E���  ����zt*���� *   3ҋEf��E������M��"����E��  �M�M�U�U��	�E����E��M�M؋U���U�}� ts�E����ti�M���%��P�U��P��&������tH�   �� �U��
��u,����� *   3ɋUf�
�E������M������E��.  �	�E����E��o����M�+M�MЋUR�EP�M�Q�URj�M��a%��� �HQ��E��}� u*���� *   3ҋEf��E������M��!����E��   �M��MȍM������E��   �   �M���$����   �����    u�MQ�������EčM�������E��j�`j j j��URj	�M��$��� �HQ��E��}� u!����� *   �E������M������E�� ��U����U��M��j����E���M��]�����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���T�E�    �} u�} t�} t�} w	�E�    ��E�   �E��E�}� u&h8�hpjj h�   h��j���������u̃}� u3�G���    j h�   h��h�h8�������   �  �} tY3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E��M���Qh�   �U��R�d������} t	�E�     �MQ�M������U;Uv�E�E���M�M�U�U��}����w	�E�   ��E�    �E�E�}� u&h�hpjj h  h��j���������u̃}� u@�-���    j h  h��h�h��x�����E�   �M������E���  �M��!��P�U�R�EP�MQ������E��}��uy�} tY3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E܋M���Qh�   �U��R�������h��� �EčM������E��G  �M����M��} �  �U�;U��   �}���   3��Mf��}�tJ�}���tA�}v;�U��9h�s
�h��E��	�M���M؋U���Rh�   �E��P�|������M�;Mw	�E�   ��E�    �UԉUЃ}� u&h<�hpjj h  h��j�(�������u̃}� u=�}��� "   j h  h��h�h<��������E�"   �M�������E��9�M�M��E�P   3ҋE��Mf�TA��} t�U�E���M̉M��M�������E���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��=4� uh��EP�MQ�UR���������j �EP�MQ�UR������]��������������������������������U��j �EP�MQ�UR�EP�MQ������]��������������U����E���E��M�M��U����U�t�E����t�U����U����}� t�E����u�E�+E������E��]������������������������U��EP�MQ�UR�EP������]��������������������U���   ���3ŉE��E�    �E�    �} t�} u3���  �} t	�E�   ��E�    �EĉEȃ}� u#ht�hpjj jfh��j��������u̃}� u.�e���    j jfh��h�ht����������M  �UR�M������} �9  �M������ �   �ჼ�    ��   �U�;Usv�E����   ~"����� *   �E������M������E���  �UU��E��
�U��E��M���M�}� u�U��U��M��P����E��  �E����E�낋M��M��M��/����E��  �|  �M��#����zt��   �} v�EP�MQ�������E�U�Rj �EP�MQ�UR�EPj �M�������QR��E��}� t3�}� u-�EE��H���u	�U����U��E��E��M������E���  ����� *   �E������M��s����E���  ��  �M�Qj �UR�EPj��MQj �M��Q����BP��E��}� t�}� u�M����M��M������E��q  �}� u����zt"�J��� *   �E������M�������E��>  �U�;U�  �E�Pj �M�������QtR�E�Pj�MQj �M������BP��E؃}� t�}� t"����� *   �E������M��x����E���  �}� |�}�v"���� *   �E������M��J����E��  �M�M�;Mv�U��U��M��)����E��~  �E�    ��EЃ��EЋM����M��U�;U�}4�EE��MЊT��EE����u�U��U��M�������E��)  벋E���E������M��M��M������E��  ��   �M������   �����    uq�E�    �M�M��	�Uԃ��UԋE����t:�U��=�   ~"���� *   �E������M��=����E��   �M̃��M�볋ỦU��M������E��t�j�E�Pj j j j��MQj �M������BP��E��}� t�}� t�'��� *   �E������M�������E���M����M��M������E���M������M�3��I�����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���4�E�    �} t�} w�} u�} t	�E�    ��E�   �E��E�}� u&h8�hpjj h@  h��j���������u̃}� u3�'���    j h@  h��h�h8��r�����   �  �} tU�U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U��E�Ph�   �M��Q�H������} t	�U�    �E;Ev�M�M���U�U�E�E��}����w	�E�   ��E�    �M�M�}� u&h�hpjj hL  h��j���������u̃}� u3����    j hL  h��h�h��h�����   �  �EP�M�Q�UR�EP�f������E��}��uf�} tT�M� �}�tH�}���t?�}v9�U��9h�s
�h��E��	�M���M܋U�Rh�   �E��P�������o��� �&  �M����M��} �  �U�;U��   �}���   �E�  �}�tI�}���t@�}v:�M��9h�s�h��U��	�E���E؋M�Qh�   �U��R�������E;E�v	�E�   ��E�    �MԉMЃ}� u&h�hpjj hd  h��j�@�������u̃}� u0���� "   j hd  h��h�h��������"   �(�E�E��E�P   �MM��A� �} t�U�E���E̋�]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�������]����������������������U��j �EP�MQ�UR�EP�MQ�������]��������������U��j�h`�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j�L������E�    �E�    �	�E���E�M�;��N  �U䡜�<� ��   �M�����H��   ��   �U䡜���Q�� �  ��   �}�~�}�}�E��P�������u��   �M����P�M�Q�R������U䡜���Q��   t�E����R�E�P�N�����0����M�����E��   �{jZh8�jj8�W������E܋M���E܉��}� tNj h�  �M������ P�������M������ P� �M�����E��M��A    ������}� tB�U��B% �  �M��A�U��B    �E��@    �M��    �U��B    �E��@�����E������   �j�������ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������U���X�E�    �$��E��E�    �E�    �E�    �} u#h��hpjj jDh��j��������u̃} u#h�hpjj jEh��j�]�������u̃} u#hl�hpjj jFh��j�4�������u̋M��� u�E���E��M��U��}�at8�}�rt�}�wt�<�E�    �E����E��   �E�  �M����M��   �E�	  �U����U��v3�t	�E�   ��E�    �M܉M؃}� u#h8�hpjj jbh��j��������u̃}� u-�����    j jbh��h��h8��& ����3���  �E�   �E���E�M����<  �}� �2  �E��M�U�� �U�}�T��  �E���xj�$�Dj��  �U���t	�E�    �'�E����E��M�����M��U��ʀ   �U��E�����E��  �M��� �  t	�E�    ��U��� �  �U��  �E�% �  t	�E�    ��M��� @  �M��u  �}� t	�E�    ��E�   �U��� @  �U��N  �}� t	�E�    ��E�   �E�%�����E��(  �}� t	�E�    ��E�   �M��� �M��  �}� t	�E�    ��E�   �U����U���   �E�%   t	�E�    ��M���   �M��   �U���@t	�E�    �	�E���@�E��   �M��ɀ   �M��   �E�   �E�    �|3�t	�E�   ��E�    �EԉEЃ}� u&h8�hpjj h�   h��j�1�������u̃}� u0����    j h�   h��h��h8��������3��  �����}� �w  �U��� u�M���M��j�URhh���������t|3�t	�E�   ��E�    �MȉMă}� u&h8�hpjj h�   h��j�y�������u̃}� u0�����    j h�   h��h��h8�������3���  �E���E�M��� u�E���E��M���=t|3�t	�E�   ��E�    �M��M��}� u&h8�hpjj h�   h��j�ӽ������u̃}� u0�(���    j h�   h��h��h8��s�����3��1  �E���E�M��� u�E���E��jhl��MQ���������u�U���U�E�   �E���   jht��MQ��������u�U���U�E�   �E��   jh���MQ�j�������u�U���U�E�   �E��|3�t	�E�   ��E�    �U��U��}� u&h8�hpjj h  h��j諼������u̃}� u0� ���    j h  h��h��h8��K�����3��	  �M��� u�E���E��M���u	�E�   ��E�    �E��E��}� u&h��hpjj h  h��j��������u̃}� u-�h���    j h  h��h��h��������3��th�  �UR�E�P�MQ�U�R�������t3��O�|����|��M�M��U��E��B�M��A    �U��    �E��@    �M��A    �U��E��B�E���]ÍI �d�d"f�ef�e�e�e�d9e`ee2f 	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������SVW�T$�D$�L$URPQQh`md�5    ���3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C������   �C賹���d�    ��_^[ËL$�A   �   t3�D$�H3������U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�I���3�3�3�3�3���U��SVWj RhnQ����_^[]�U�l$RQ�t$������]� ����������������������������������������������������������������������������������������������U��H  ������3ŉE��} tǅ����   �
ǅ����    ������������������ u#h��hpjj j\hȪj辶������u̃����� u.�����    j j\hȪh8�h���^���������  �U������������P��������������������y }�������B    jj ������P�*����������������� }����  ��������������������P��L$�����������������B%  u������������+A�Y  �������������
+H�������������B����  ���������_  ��������������������P��|0 �8  �������������
+H�鉍�����������z u��������  �  j ��������������������P��D
,P�L
(Q������R��������������������������������������P�������������������������������;T(u������������������;T,t����!  j ������Ph   ������Q��������������������P��R����u�����  j ������P������Q�.�������}����  ������;�����v����  �������������������������������������������� ��   ������������9�����ss���������u5������������9�����s�������H��
u������������������������X���������������������������P���������������+ʋ�3�������������  ��������������������P��T��   tO�������H���������������������������������;s���������
u�����������������#�������B%�   u�����    ����$  ������ u�������  �������Q����  �������x uǅ����    �  �������������+B������A��������������������������P��T��   �^  jj ������P�������;�������   �������Q������������������H���������������������������;�����s���������
u���������������ċ������Q��    t���������������   j ������Q������R�D�������}�����   ������   w*�������H��t�������B%   uǅ����   ��������Q��������������������������P��D
��t����������������������u�������艅����������+�������������������u�������艅����������������M�3��9�����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h�hpjj j0hȪj�=�������u̃}� u+�����    j j0hȪh(�h������������@�UR�F������E�    �EP�w������E��E������   ��MQ� �����ËE܋M�d�    Y_^[��]������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u�~����     ����� 	   �����  �} |�E;\�s	�E�   ��E�    �M��M܃}� u#h`hpjj jAh`�j�ά������u̃}� u9�
����     ����� 	   j jAh`�h��h`�f���������L  �E���M������P��D
��t	�E�   ��E�    �M؉Mԃ}� u#h�`hpjj jBh`�j�0�������u̃}� u9�l����     �z���� 	   j jBh`�h��h�`�����������   �EP�%������E�    �M���U������P��L��t�UR�EP�MQ�(������E��D� ���� 	   �ܰ���     �E�����3�u#h(ahpjj jMh`�j�a�������u��E������   ��MQ�������ËE�M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������U����EP�c������E��}��u:������ 	   3�u#hЫhpjj jkh`�j�L�������u̃����   �E�    �E�    j�E�P�M�Q�U�R�E�P����u��P�Ϩ��������   �E��E�U��MQ�U�R�E�P�M�Q�U�R����u��P萨��������g�}� t&j j �E�P�M�Q�U�R�������    ����;�E���M������P��D
����M���U������P��D�E��]������������������������������������������������������������������������������������U���X�E�    �$��E��E�    �E�    �E�    �} u#h��hpjj jDh��j趨������u̃} u#h�hpjj jEh��j荨������u̃} u#hl�hpjj jFh��j�d�������u̋M��� u�E���E��M��U��}�at8�}�rt�}�wt�<�E�    �E����E��   �E�  �M����M��   �E�	  �U����U��v3�t	�E�   ��E�    �M܉M؃}� u#h8�hpjj jbh��j貧������u̃}� u-�����    j jbh��h\�h8��U�����3���  �E�   �E���E�M����<  �}� �2  �E��M�U�� �U�}�T��  �E���H��$����  �U���t	�E�    �'�E����E��M�����M��U��ʀ   �U��E�����E��  �M��� �  t	�E�    ��U��� �  �U��  �E�% �  t	�E�    ��M��� @  �M��u  �}� t	�E�    ��E�   �U��� @  �U��N  �}� t	�E�    ��E�   �E�%�����E��(  �}� t	�E�    ��E�   �M��� �M��  �}� t	�E�    ��E�   �U����U���   �E�%   t	�E�    ��M���   �M��   �U���@t	�E�    �	�E���@�E��   �M��ɀ   �M��   �E�   �E�    �|3�t	�E�   ��E�    �EԉEЃ}� u&h8�hpjj h�   h��j�`�������u̃}� u0�����    j h�   h��h\�h8�� �����3��  �����}� �w  �U��� u�M���M��j�URh��]�������t|3�t	�E�   ��E�    �MȉMă}� u&h8�hpjj h�   h��j訤������u̃}� u0������    j h�   h��h\�h8��H�����3���  �E���E�M��� u�E���E��M���=t|3�t	�E�   ��E�    �M��M��}� u&h8�hpjj h�   h��j��������u̃}� u0�W����    j h�   h��h\�h8�������3��1  �E���E�M��� u�E���E��jh ��MQ���������u�U��
�U�E�   �E���   jh,��MQ���������u�U���U�E�   �E��   jh@��MQ��������u�U���U�E�   �E��|3�t	�E�   ��E�    �U��U��}� u&h8�hpjj h  h��j�ڢ������u̃}� u0�/����    j h  h��h\�h8��z�����3��	  �M��� u�E���E��M���u	�E�   ��E�    �E��E��}� u&h��hpjj h  h��j�B�������u̃}� u-�����    j h  h��h\�h���������3��th�  �UR�E�P�MQ�U�R���������t3��O�|����|��M�M��U��E��B�M��A    �U��    �E��@    �M��A    �U��E��B�E���]Ë�~�~���{W��~
1�~� 	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U������]��E�E��M������U�ҁ�   �ʉM��E���]����������������U������]��E�E��M��M�U��%����M���ҁ�   �M��E���]���������������������U������]��E�E��M������U��   �ʉM��E���]������������������U������]��E�E��M�M�U��U��E��������U�%   �ȋU��
�E���]�����������������U���E%�  =�  u3���   ]�������������������U����E%�  =�  uP���E�$�\������E��}�t�}�t�}�t��   �   �   �   �   �   �   �   �M�� �  �M��U���  u+�E����u�} t�}� t	�E�   ��E�   �E��B�E��������Dz�}� t	�E�    ��E�@   �E���}� t	�E�   ��E�   �E��]�����������������������������������������������������������������U���E%�  =�  u�M����u�} u�U���  ���  u�   �3�]�����������������U������]�h��  h?  ��������E��E%�  =�  ��   ���E�$�������E��}� ~C�}�~�}�t�5h��  �M�Q�������E�   �U�R���E�$j%��������   �E�P�E��s���$���E�$j%j螚�����q�E��������Dz)�M�Q�p������$���E�$j%j�g������:�U�R���E�$�����؃��E���E��E��]�h��  �M�Q��������E��]���������������������������������������������������������������������������������U���$���]�h��  h?  �u������E��E%�  =�  t�M���  ���  ��   �U���  ���  u�E����u(�} u"�M���  ���  uC�U����u�} t3�E�P�E�E���$���E�$���E�$j&j�3�����$�\  �M���  ���  t�U���  ���  u%�E�P���E�$���E�$j&�������  �E�E������Dzh��  �M�Q�l������E��  �E��������Dz$�E�   �E�]����z	�E�    ��E�   ����]����z�E�]����At���]����Au-�E�]����z �U���U�E�E��} u	�M����M��P���]����z�E�]����{���]����Au+�E�]����Au�U���U�E�E��}� u	�M����M��U���  uv�E�����u�}� tf�M�Q���E��$��������]�U���   R���E��$�ڱ�����]�E�P���E��$���E�$���E�$j&j�l�����$�   �}�  �u�}� t�}�  ��ui�}� uc�M�Q���E��$�Y������]܋U��   R���E��$�V������]�E�P���E��$���E�$���E�$j&j������$�h��  �M�Q�|������E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EP���E�$������]�������U��EPj �MQh�]������]���������������������U���0�E�    3��EԉE؉E܉E��E�E�E�MЉM��} t	�E�   ��E�    �U��U�}� u&h��hpjj h�  hȎj��������u̃}� u.�\����    j h�  hȎh��h������������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]��������������������������������������������������������������������U��EP�MQ�URh�]�F�����]�������������������U��EPj �MQhsa������]���������������������U��EP�MQ�URhsa�������]�������������������U���@�E�    3��EĉEȉẺEЉEԉE؉E܍M��M��} t	�E�   ��E�    �U��U�}� u#h��hpjj jphȎj�J�������u̃}� u.�����    j jphȎhx�h�������������  �} t	�E�   ��E�    �M��M�}� u#hX�hpjj juhȎj�ѓ������u̃}� u.�&����    j juhȎhx�hX��t���������   �E��@����M��AB   �U��E�B�M��U��EP�MQ�UR�E�P�w������E�} u�E��Q�M��Q���U�E��M�H�}� |"�U���  3Ɂ��   �M��U�����M����U�Rj �S������E��E��]���������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR������]����������������������U����EPj �MQ�UR�EPh�]�/������E��}� }	�E�������M��M��E���]�����������������������������U����EP�MQ�UR�EP�MQh�]�ͳ�����E��}� }	�E�������U��U��E���]���������������������������U���@�E�    3��EĉEȉẺEЉEԉE؉E܍M��M��} t	�E�   ��E�    �U�U��}� u#h��hpjj jphȎj�*�������u̃}� u.�����    j jphȎh��h�������������W  �} t�} u	�E�    ��E�   �M�M�}� u#hP�hpjj jshȎj諐������u̃}� u.� ����    j jshȎh��hP��N����������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R�U���E��} u�E��{�}� |X�E��H���M�U��E�B�}� |!�M��� 3�%�   �E��M�����E����M�Qj �������E��}��t�E���UU�B� �E��x }�����������]�����������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP�MQ�E�����]��������������U���0�E������E�    �} t	�E�   ��E�    �E�E��}� u&h�hpjj h  hȎj荎������u̃}� u1������    j h  hȎhȭh��-���������'  �} u�} u�} u3��  �} t�} v	�E�   ��E�    �U�U�}� u&h8�hpjj h  hȎj��������u̃}� u1�D����    j h  hȎhȭh8�����������  �M;M��   ������U��EP�MQ�UR�E��P�MQh``�y������E��}��u~�}�t\�}���tS�U��;UsH�E���M+�9h�s�h��U���E���M+ȉM�U�Rh�   �E�M�TR�������n����8"u
�d����M�������  �`�P�����U��EP�MQ�UR�EP�MQh``�Ů�����E��UU�B� �}��u"�}�u�����8"u
�����M������f  �}� ��   �   k� �M� �}�tH�}���t?�}v9�U��9h�s
�h��E��	�M���M��U�Rh�   �E��P�8������}��uz3�t	�E�   ��E�    �U܉U؃}� u&h��hpjj hB  hȎj��������u̃}� u.�7���� "   j hB  hȎhȭh����������������z�}�t\�}���tS�M���;MsH�U����E+�9h�s�h��M���U����E+EԋM�Qh�   �U��E�LQ�Q������}� }	�E�������U��UЋEЋ�]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EPj �MQ�UR�EPhsa�������E��}� }	�E�������M��M��E���]�����������������������������U����EP�MQ�UR�EP�MQhsa譫�����E��}� }	�E�������U��U��E���]���������������������������U���$�E������} t	�E�   ��E�    �E��E�}� u&h�hpjj h�   hȎj�$�������u̃}� u1�y����    j h�   hȎh�h�������������  �} t�} v	�E�   ��E�    �U��U�}� u&h8�hpjj h�   hȎj蟈������u̃}� u1������    j h�   hȎh�h8��?���������s  �MQ�UR�EP�MQ�URh``�B������E��}� }^�   k� �U�
 �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U�E�Ph�   �M��Q�������}��uz3�t	�E�   ��E�    �E�E��}� u&h��hpjj h�   hȎj蔇������u̃}� u.������ "   j h�   hȎh�h���4���������k�}� |b�}�t\�}���tS�U���;UsH�E����M+�9h�s�h��U���E����M+ȉM܋U�Rh�   �E��M�TR�������E���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP�*�����]������������������U���8  ���3ŉE�ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    �EP�� ����b���ǅ����    �������d����} tǅ���   �
ǅ���    �������$�����$��� u&h�hpjj h  hx�j�1�������u̃�$��� uI�����    j h  hx�hخh��������ǅ���������� ���������������W  �E��\�����\����Q��@��   ��\���P�������������������t-�������t$�������������������P�������
ǅ����������H$�����х�uV�������t-�������t$�������������������P���0����
ǅ0������0����B$�� ���ȅ�tǅ,���    �
ǅ,���   ��,�����P�����P��� u&hh�hpjj h	  hx�j贃������u̃�P��� uI�����    j h	  hx�hخhh��Q�����ǅ���������� ���聝����������  �} tǅ���   �
ǅ���    �������H�����H��� u&h��hpjj h  hx�j��������u̃�H��� uI�]����    j h  hx�hخh��������ǅ���������� ����؜���������1  ǅ����    ǅ����    ǅ����    ǅ����    ǅ|���    �E��������������������E���E������ ��  ������ ��  �������� |%��������x�������������(����
ǅ(���    ��(�����������������������������������������@�����@����%  ��@����$�0�ǅ����    �� ��������P������R�����������   ������P�MQ������R�3  ���E��������U���U��������tǅ���   �
ǅ���    �������8�����8��� u&h�hpjj h�  hx�j�	�������u̃�8��� uI�[����    j h�  hx�hخh�覿����ǅ���������� ����֚���������/  ������P�MQ������R�V  ����  ǅ����    ������������������������������������ǅ����    ǅ��������ǅ����    �  �������������������� ������������wj��������h��$�P����������������E���������������4���������������#�������ɀ   ����������������������  ��������*u:�MQ�x����������������� }���������������������؉������k�����
�������DЉ������  ǅ����    �  ��������*u'�UR������������������ }
ǅ���������k�����
�������TЉ������F  ��������������������I������������.�3  �����������$�|��M���lu�E���E��������   �����������������������   �E���6u,�U�B��4u �M���M�������� �  �������   �E���3u)�U�B��2u�M���M������������������S�E���dt7�U���it,�M���ot!�E���ut�U���xt�M���Xu�ǅ����    ������#�������� ���������������   ��������  ��������������������A������������7�)
  �����������$���������%0  u��������   ��������������  t[ǅ ���    �EP�O�����f��`�����`���Qh   ������R������P�y������� ����� ��� t
ǅ����   �2�MQ蜓����f��x����   k� ��x���������ǅ����   �������������J	  �EP�Y����������������� t�������y u#�p�������������P�e������������e��������   t/�������B��������������+���������ǅ����   �(ǅ����    �������B��������������������  ������%0  u��������   �������������uǅX���������������X�����X����������MQ�Y�������������������  ��   ������ u�t�������ǅ����   �������������������������������������������� t���������t��������������뾋�����+��������������u������ u�p��������������������������������������������������� t���������t��������������뾋�����+������������*  �MQ�9�������D�����������   3�tǅT���   �
ǅT���    ��T�����L�����L��� u&h�hpjj h�  hx�j��y������u̃�L��� uI�E����    j h�  hx�hخh�萸����ǅ���������� ���������������	  �_  �������� t��D���f������f����D����������ǅ����   �%  ǅ����   �������� ��������������@������������������ǅ|���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Zh�  hp�j��������]  R�t���������������� t ��������������������]  ��|����
ǅ�����   �U���U�E�H��P��������������� ����e���P������P������Q������R��|���P������Q������R�   k���0�R��Ѓ�������%�   t6������ u-�� ��������P������Q�   k�	��0�Q��Ѓ���������gu:������%�   u-�� �������P������Q�   ����0�P��Ѓ����������-u ������   ��������������������������R�\�������������  ��������@������ǅ����
   �   ǅ����
   �   ǅ����   ǅ����   �
ǅ����'   ǅ����   ��������   t2�   k� Ƅ����0��������Q�   �� ������ǅ����   �)ǅ����   ������%�   t��������   �������������� �  t�EP�f������������������   ��������   t�UR�;������������������   �������� tE��������@t�UR�Ռ��������������������EP蹌��������������������@��������@t�UR萌�������������������EP�u�����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ������������������ }ǅ����   �%���������������������   ~
ǅ����   �����������u
ǅ����    �   i��  �������������������������������������������� �������������   �������RP������R������P�č����0�������������RP������Q������R� ���������������������9~���������������������������������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0�������������������� �b  ��������@tv��������   t�   k� Ƅ����-ǅ����   �L��������t�   k� Ƅ����+ǅ����   �%��������t�   k� Ƅ���� ǅ����   ������+�����+�������l�����������u������Q�UR��l���Pj ��	  ����d���Q������R�EP������Q������R�"
  ����������t'��������u������R�EP��l���Qj0�	  �������� ��   ������ ��   ǅ<���    ��������t�����������h�����h�����������h�������h��������� ��   ��t���f�f��r�����r���Rj�E�P��4���Q��������<�����t�������t�����<��� u	��4��� uǅ���������*��d���P������Q�UR��4���P�M�Q�	  ���N����(��d���R������P�MQ������R������P��  �������� |'��������t������R�EP��l���Qj �X  �������� tj������R�T����ǅ����    ������������������ ���袊���������M�3��B�����]Ð��c���Z�i������ϥ������ �I 2������ �G�W�֩��"�a�v�x�B����������l�   	
������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E����U�
�E��A��Q�]��������������������U��E����U�
�E��A�]�������U��E����U�
�E�f�A�]����������������������U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�������E��}��u�M�������U����M���]�������������������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��|�U�    �E�E��M���M�}� ~N�U��E��MQ�UR�E�P�w������M���M�U�:�u�E�8*u�MQ�URj?�L�������띋E�8 u�M�U���]������������������������������������������������U��� �=4� ��  �} t	�E�   ��E�    �E�E��}� u#hԸhpjj jXh��j��f������u̃}� u0�F����    j jXh��h �hԸ蔥���������/  �} t	�E�   ��E�    �U�U�}� u#hp�hpjj jYh��j�vf������u̃}� u0�ˬ���    j jYh��h �hp������������   �M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���M�U���U�E���t�M��U�;��l����E��M�+���j �UR�EP蕒������]��������������������������������������������������������������������������������������������������������������������������������U���@�EP�M��n���} t	�E�   ��E�    �M��M�}� u#hԸhpjj j4h��j�d������u̃}� u=�����    j j4h��h�hԸ�U������E�����M��~���E���  �} t	�E�   ��E�    �E�E�}� u#hp�hpjj j5h��j�*d������u̃}� u=�����    j j5h��h�hp��͢�����E�����M��~���E��;  �M��������   �����    ��   �M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���M�U���U�E���t�M��U�;��l����n�Ef�f�M��M��=���P�U�R�U`����f�E��E���E�Mf�f�U�M�����P�E�P�(`����f�E��M���M�U���t�E��M�;�t��U��E�+ЉUЍM���|���EЋ�]����������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h �h�Ld�    P��SVW���1E�3�P�E�d�    �=<� uEj�b�����E�    �=<� u�(  �<����<��E������   �j�ٚ����ËM�d�    Y_^[��]�������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j��a�����E�    �EP�_   ���E��E������   �j�'�����ËE�M�d�    Y_^[��]��������������������������������������������U����E�    j h9  h8�h��h���E�P��e����P�7k�����}� u3��  �M�Q;|�u�E�H;����  �=@� �G  �����uO���P���Q���R���Pj ���Q���R���P�M�QRjj�i  ��,�G���P���Q���R���P���Qj j ���R�E�HQj j�   ��,�����uO���P���Q���R���Pj ���Q���R���P�M�QRjj ��
  ��,�G���P���Q���R���P���Qj j ���R�E�HQj j �
  ��,�   �E�   �E�   �E�   �E�   �U�zk}�E�   �E�   �E�
   �E�   j j j jj j �E�P�M�Q�U�BPjj�
  ��,j j j jj j �M�Q�U�R�E�HQjj ��	  ��,���;��}K�E�H;��|�U�B;��~3���   �M�Q;��~�E�H;��}
�   �   �F�U�B;��|�M�Q;��~
�   �   �E�H;��~�U�B;��}3��a�MkQ<�E�ʋUiB  �i��  �M�U�B;��u�M�;��|	�   ��3����U�;��}	�   ��3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����z���M�]������������������U��萑���M�]������������������U�������M�]������������������U��j�h��h�Ld�    P��SVW���1E�3�P�E�d�    j��\�����E�    �J   �E������   �j������ËM�d�    Y_^[��]��������������������������������U��j�h �h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    j�\�����E�    �|����E�j h�   h8�h��h���E�P�b����P�e����j h�   h8�h��h���M�Q�M`����P�e����j h�   h8�h��h0��U�R�~����P�de�����<����E��@�    �����������|�hh��~|�����E�}� t�M������  �=8� tj�8�P��h�����8�    hH��@����=  �@�   kH�<�M������tk��<E��E������t$�=�� t�E�   ���+��k�<�E���E�    �E�    �M�Qj j?�   k� �M܋Rj�hL�j �E�P���t"�}� u�   k� �   k�?�E܋� ��   k� �   k� �U܋
� �U�Rj j?�   �� �M܋Rj�h��j �E�P���t"�}� u�   �� �   k�?�U܋
� ��   �� �   k� �E܋� �E�   ��   �=8� t"�8�P�M�Q��������u�E�   �   �=8� tj�8�R�g����h  hl�j�E�P臂������P�cT�����8��=8� u	�E�   �Aj h   h8�h��h���M�Q�U�R�>�������P�8�P襟����P��b�����M�Q�ӧ�����U�R�ɖ�����E�P�ч�����E������   �j������Ã}� ��  j h3  h8�h��h��j�M�Qj@�   k� �M܋R虣����P�Tb�����E���E�M����-u�Eȃ��EȋM���M�U�R�Ӝ����i�  �E��M����+t�E����0|�U����9�M���M��ԋU����:��   �M���M�U�R�z�����k�<E��E��M����0|�E����9�U���U��ߋE����:u<�U���U�E�P�0�����E��E��M����0|�E����9�U���U��߃}� t�E��؉E��M����t	�E�   ��E�    �}� t@j hj  h8�h��hH�j�E�Pj@�   �� �U܋
P�1�����P��`������   �� �U܋
�  �M�Q�ӥ�����U�R�ɔ�����M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���VW�E�    �}�K  �E%  �yH���@��u�E��d   ����u#�El  ���  ����t�U�����E���M�����U�E���E��M��Fi�m  M��E���������E����d   ��+��E+  ���  ����D1�   ���U��U�;U�E+E��M��k�U�ЉU���E+E�kMM�ȉM��}ud�U��  �yJ���B��u�E��d   ����u#�El  ���  ����t�U�����E���M�����U��E�;E�~	�M����M��b�U��  �yJ���B��u�E��d   ����u#�El  ���  ����t�U�����E���M�����U�E�E��M�M �M��}u2�U����kE$<E(k�<M,i��  U0����E�|��   �M����kU$<U(k�<E,i��  M0���j h�  h8�h��h0��U�R�u����P��\����iE��  �����y#����� \&������������*�=�� \&|���- \&������������U���_^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U�츜�]�������U�츠�]�������U�츘�]�������U��(�]�������U����} t	�E�   ��E�    �E��E��}� u#h�hpjj j$hP�j�nP������u̃}� u-�Ö���    j j$hP�h��h��������   ��U����3���]���������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u#hسhpjj j-hP�j�O������u̃}� u-�����    j j-hP�h(�hس�Q������   ��U����3���]���������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u#hH�hpjj j6hP�j��N������u̃}� u-�C����    j j6hP�hx�hH�葍�����   ��U����3���]���������������������������������������������������U����} t�} w�} u�} t	�E�    ��E�   �E��E��}� u#h��hpjj j?hP�j�N������u̃}� u0�q����    j j?hP�h`�h��迌�����   �_  �} t�   k� �M� �} t	�E�   ��E�    �U�U��}� u#h|�hpjj jDhP�j�M������u̃}� u0�����    j jDhP�h`�h|��/������   ��   �} t�}t	�E�    ��E�   �M�M�}� u#h��hpjj jEhP�j�M������u̃}� u-�`����    j jEhP�h`�h��讋�����   �Q�E��(�Q��v�������U��} u3��,�E�;Mv�"   ��U��(�P�MQ�UR� �������]�������������������������������������������������������������������������������������������������������������������������������������������U��Qh  �EP��������u�M��_t	�E�    ��E�   �E���]�����������������������U��Qh  �EP�ˀ������u�M��_t	�E�    ��E�   �E���]�����������������������U����EP�M��U���M��\�����U���   �P�� �  �M��M��2e���E���]�������������������������������U��h  �EP������]����������U��h  �EP������]����������U��Q�E��	u	�E�@   �j@�MQ�������E��E���]������������������U��j �EP�����]�������������U��Qh  �EP�{������u�M��_t	�E�    ��E�   �E���]�����������������������U��Qh  �EP�+������u�M��_t	�E�    ��E�   �E���]�����������������������U��j�EP��~����]�������������U��h  �EP�~����]����������U��j�EP�~����]�������������U��hW  �EP�|~����]����������U��j�EP�_~����]�������������U��j�EP�?~����]�������������U��j�EP�~����]�������������U��h�   �EP��}����]����������U��j �EP������]��������������U��h  �EP�}����]����������U��h  �EP�}����]����������U��Q�E=�   s	�E�   ��E�    �E���]�����������U��Q�E��	u	�E�@   �j@�MQ�<}�����E��E���]������������������U��j �EP�}����]�������������U��j�EP��|����]�������������U��h  �EP��|����]����������U��j�EP�|����]�������������U��hW  �EP�|����]����������U��j�EP�o|����]�������������U��j�EP�O|����]�������������U��j�EP�/|����]�������������U��h�   �EP�|����]����������U��Q�E�    ��E����E��M���M�U�;Us�E���t�ڋE���]�����������������������U���  ���3ŉE��= � t3��M�3��e����]�� ��X  ����   Vh����5���tjh  ������QP�(��tSh  ������P������P��  ����t4h 	  j ������P�օ���   ����Wujj ������P�օ�ugh 
  j h`��օ�uU����WuHh  ������Pj �(��t0h  ������P������P�C  ����tjj ������P�օ�u3�^�M�3��d����]�������������������������������������������������������������������������������������������U���$  ���3ŉE�S��Wh   j hX��Ӌ���u,����WuWWhX��Ӌ���u_3�[�M�3��Vc����]�V�5�hx�W�։�������tJh��W�։�������t8h��W�։�������t&������Pjj h��h  ���������tW�H^_3�[�M�3���b����]Í�����ǅ����  P������P������Pj h ���������������������������W�H��u�������u���������u����r�If9�M�����x���f��M����\t�\   f��M����A���+����Q����A=  �C�������M��������M��������M��������M �������M���� ���M����$���M����(���M���f�,�h 	  f��M���������j P�Ӌ���u����WujV������P�Ӌ��M���^_3�[�a����]������������������������������������������������������������������������������������������������������������������������������������������������������U���  ���3ŉE��E������V�uh   Qh   ������Qh   ������Qj�M�QP��d����$��t3�^�M�3��`����]�hH�������j	P��������u�h<�������jP�ш������u�������P������P������P�E�P�uV�"U���M������3�@^�"`����]������������������������������������������������������������������U��E��D3��     �ES�]jf�K�E�PS�D��u3�[��]��u�u�u��(��t�M��MZ  f9uًA<��~ҁ<PE  V�4t^3�[��]��F+��V��$�3�W3���t�;�r	��+�;X�rG��(;�r�;�t]G�=!� u �=� uJ���������t<�!����hx�P����t�M�Qj j �M�Qj j j �u�Ѓ� ��u	_^3�[��]ËM�3ۉ]��=A�2�}  �M��U�Rh`�S��P���c  �M�U�SSS�RVW�P ���B  �M�U��]�R��@h�Є��!  �M����  ��P����   �M��U�j R�U��R�UR�@�U�Rj �Є���   �E;�u�M�;�w	�E��;�r�M���P��u��   �E�����   =�����   ��Pj �(P�$�؅��}   �M��U�SRj ��U�j j R�@�Є�tP+u�;3rI�M��   ;�v
;4�r@;�r��D���U�M%��� j j j ��M�R�u��u܋@p�Є�t�E�   Sj �(P��M����]�M��P@�M��R8�M���R,_^��[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���<�} t�} v	�E�   ��E�    �E�E��}� u#hhhpjj jh��j�h=������u̃}� u0轃���    j jh��h�hh�|�����   �  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R��c�����} t	�E�   ��E�    �E�E�}� u#h�^hpjj jh��j�<������u̃}� u0�߂���    j jh��h�h�^�-{�����   �  �U�U��E�E��}� v�M����t�E����E��M����M��܃}� ��   3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E��M���Qh�   �U��R��b��������t3�t	�E�   ��E�    �U܉U؃}� u#hP�hpjj j h��j�u;������u̃}� u0�ʁ���    j j h��h�hP��z�����   �  �M��Uf�f��M���UċE����E��M���M�}� t�U����U�t�ƃ}� ��   3��Mf��}�tJ�}���tA�}v;�U��9h�s
�h��E��	�M���MԋU���Rh�   �E��P�a����� _��t3�t	�E�   ��E�    �EЉẼ}� u#hP_hpjj j*h��j�W:������u̃}� u-謀��� "   j j*h��h�hP_��x�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9h�s�h��U���E+E����M+ȉMȋU���Rh�   �E+E��M�TAR�`����3���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���8�} u�} u�} u3��  �} t�} v	�E�   ��E�    �E�E��}� u#hhhpjj jh��j�?8������u̃}� u0�~���    j jh��h�hh��v�����   �  �} u`3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R�^����3��&  �} ��   3��Mf��}�tJ�}���tA�}v;�U��9h�s
�h��E��	�M���M�U���Rh�   �E��P�K^�����} t	�E�   ��E�    �M�M��}� u#h�^hpjj jh��j��6������u̃}� u0�Q}���    j jh��h�h�^�u�����   �I  �E�E��M�M��}�u?�U��Ef�f�
�U���E̋M����M��U���U�}� t�E����E�t���   ��k����t+�M;Mr#h _hpjj j+h��j�A6������u̋E��Mf�f��E���MȋU����U��E���E�}� t�M����M�t�U���Ut뻃} u3��M�f��}� ��   �}�u3ҋE�Mf�TA��P   �J  3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E܋M���Qh�   �U��R�x\����� _��t3�t	�E�   ��E�    �U؉Uԃ}� u#hP_hpjj j>h��j�"5������u̃}� u-�w{��� "   j j>h��h�hP_��s�����"   �r�}�tj�}���ta�M+M���;MsS�U+U����E+�9h�s�h��M���U+U����E+EЋM���Qh�   �U+U��E�LPQ�[����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E���]����U����E�    �E�E��}� |,�}�~�}�t��$��M��U�$��~�$��E��t3�t	�E�   ��E�    �U�U��}� u#h,�hpjj j?hp�j��2������u̃}� u+�&y���    j j?hp�hйh,��tq���������E���]�������������������������������������������������U���8�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E��}� u#h^hpjj jh��j��1������u̃}� u0�Tx���    j jh��h��h^�p�����   �v  �} u\�U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U�E�Ph�   �M��Q�xX����3��  �} ��   �U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U�E�Ph�   �M��Q�X�����} t	�E�   ��E�    �U�U��}� u#h�^hpjj jh��j��0������u̃}� u0�w���    j jh��h��h�^�fo�����   �:  �M�M��U�U��}�u=�E��M���E���M̋U����U��E���E�}� t�M����M�t���   �e����t+�U;Ur#h _hpjj j+h��j�
0������u̋M��U���M���UȋE����E��M���M�}� t�U����U�t�E���Et뽃} u�M�� �}� ��   �}�u�UU�B� �P   �D  �E�  �}�tI�}���t@�}v:�M��9h�s�h��U��	�E���E܋M�Qh�   �U��R�LV����� _��t3�t	�E�   ��E�    �U؉Uԃ}� u#hP_hpjj j>h��j��.������u̃}� u-�Ku��� "   j j>h��h��hP_�m�����"   �p�}�th�}���t_�M+M���;MsQ�U+U����E+�9h�s�h��M���U+U����E+EЋM�Qh�   �U+U��E�LQ�_U����3���]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    �E��Q�U�j j �EP�MQ�+�����E��}� u3���   �}� ~W3�uS�����3��u���rD�E���P�L9������t#h��  �M��T	R�W����P�n�����E���E�    �E��E���E�    �M�M��}� u3��u�U�R�E�P�MQ�UR�x*������u�H�F�} uj j j j j��E�Pj �M�Q��E��!j j �UR�EPj��M�Qj �U�R��E�E�P��C�����E��]����������������������������������������������������������������������������������������U����EP�M��|5���MQ�UR�EP�MQ�M��x��P�P������E��M��E���E���]����������������������������U����E�MH<�M��E�    �U��B�M��T�U���E���E�M���(�M��U��B9E�s#�M��U;Qr�E��H�U�J9Ms�E���3���]������������������������������U��j�h@�h�Ld�    P���SVW���1E�3�P�E�d�    �e��E�   �E�    �E�P�Z������u�E�    �E������E��   �M+M�MЋU�R�E�P��V�����E��}� u�E�    �E������E��}�M��Q$��   �u	�E�   ��E�    �E܉E��E������E��M�E������D�M���Eā}�  �u	�E�   ��E�    �E�Ëe��E�    �E������E���E������M�d�    Y_^[��]��������������������������������������������������������������������������������������U����E�E��M����MZ  t3��;�E��M�H<�M��U��:PE  t3�� �E����E�M����  t3���   ��]������������������������������������U��E�(�]����U���(V�(�P��E��} t	�E�   ��E�    �M�M��}� u#h�hpjj j>hH�j�n(������u̃}� u0��n���    j j>hH�h��h��g�����   ��  �E�     �}� ��  h   j hX����E��}� u����Wuj j hX����E��}� uy3�t	�E�   ��E�    �U�U�}� u#h��hpjj jVhH�j�'������u̃}� u0��m���    j jVhH�h��h���Gf�����   ��   h,��M�Q���E��}� ��   3�t	�E�   ��E�    �E�E��}� u#h��hpjj j\hH�j�'������u̃}� uD��P��X�������Sm���0j j\hH�h��h���e������P�X�����T�U�R��E�j ��E؋Eܹ(��;E�t
�U�R�Hj�EP�U���u��l���    ��l��� �3�^��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�} t,�}t&h�hpjj h�   hH�j�%������u̋M�M��} tG�U��B%   t:�M�Q��h�����U��B%�����M��A�U��B    �E��     �M��A    ��]������������������������������������U����} u#hl�hpjj j?hH�j��$������u̋M�M��U�R�:X����P�d������u3��  �\���    �� �9E�u	�E�    �#�\���    ���9E�u	�E�   �3���   �|����|��M��Q��  t3��   �E��<�,� u\j[h��jh   �G �����E�M��U��,��}� u0�E����E��M��U��Q�E��M���U��B   �E��@   �/�M��U���,��A�M��U��B��M��A   �U��B   �E��H��  �U��J�   ��]�������������������������������������������������������������������������������������������������������U��3�]����������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E���M�����P��M��E�   �U�z uXj
��#�����E�    �E�x u%j h�  �M��Q�+Q�����U�B���M�A�E������   �j
��[����Ã}� t!�U���E������P��TR� �E��M�d�    Y_^[��]��������������������������������������������������������������������U��j�h`�h�Ld�    P���SVW���1E�3�P�E�d�    �E������E�    j�l������u����:  j�"�����E�    �E�    �	�E����E��}�@��  �M��<�P� �  �U���P��E��	�M��@�M�U���P�   9E���   �M��Q����   �E�x uXj
�"�����E�   �M�y u%j h�  �U��R�yO�����E�H���U�J�E�    �   �j
�$Z����Ã}� u+�E��P� �M��Q��t�E��P��=����}� u-�M��A�U�������E����M��U�+�P���E�������}��t��   ��   h�   h�jj@j �8�����E�}� ��   �E��M��P��\��� �\��	�E��@�E�M���P���   9U�s#�E��@ �M�������U��B
�E��@    뿋M����M܋U����E܃�����P��D�U�R��j������u�E������������E������   �j��X����ËE܋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�} ��   �E;\���   �M���U������P��L����   �U���E������P��<�th�=��u<�U�U��}� t�}�t�}�t�"j j��L�j j��L�
j j��L�E���M������P��
����3����Od��� 	   �+#���     �����]���������������������������������������������������������������U����}�u��"���     ��c��� 	   ����O  �} |�E;\�s	�E�   ��E�    �M��M��}� u&h`hpjj h5  hP�j�������u̃}� u<�X"���     �fc��� 	   j h5  hP�h��h`�[��������   �E���M������P��D
��t	�E�   ��E�    �M�M��}� u&h�`hpjj h6  hP�j�x������u̃}� u9�!���     ��b��� 	   j h6  hP�h��h�`�[���������E���M������P��
��]����������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E� �E��t
�M�� �M�U�� @  t�E��   �E�M��   t
�U���U�EP���E܃}� u��P����������q  �}�u�M��@�M���}�u
�U���U��6���E��}��u�Aa���    � ���     ����#  �E�    �EP�M�Q�1:�����U���U�E����M�������P��E�D
�M����U�������P��L$�ဋU����E�������P��L$�E����M�������P��D
$$�M����U�������P��D$�E�   �E������   �K�}� u8�U����E�������P��T����E����M�������P��T�M�Q�o����Ã}� t�U��U���E������EԋM�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������U��Q�} ��   �E;\���   �M���U������P��<�um�=��uB�M�M��}� t�}�t�}�t�(�URj��L��EPj��L��MQj��L�U���E������P��U�3����^��� 	   ����     �����]��������������������������������������������������������������U��E���M������P��D
P�]�����������U����}�u�(^��� 	   3��   �} |�E;\�s	�E�   ��E�    �M��M��}� u#h`hpjj j(hؼj�k������u̃}� u*��]��� 	   j j(hؼh8�h`�V����3���E���M������P��D
��@��]�������������������������������������������������U���,�} t�} u3��  �E���u�} t3ҋEf�3���  �MQ�M��j ���M��c����ztt3�M��c��� �xtt#hP�hpjj jGhP�j�b������u̍M��wc����   �����    u*�} t�Mf��Ef��E�   �M��90���E��c  �M��2c��P�M�R�Bd��������   �M��c��� �xt~\�M��c����U;Qt|J�} t	�E�   ��E�    �E�P�MQ�M���b����BtP�MQj	�M��b����BP���u?�M��b����U;Qtr�E�H��u"��[��� *   �E������M��n/���E��   �M��gb����Bt�E�M��N/���E��{�q�} t	�E�   ��E�    �M�Q�URj�EPj	�M��"b����QR���u�P[��� *   �E������M���.���E���E�   �M���.���E���M���.����]����������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�MX����]����������������������U��j�hОh�Ld�    P���SVW���1E�3�P�E�d�    3�f�E�j������E�    �MQ�Y����f�E��E������   �j��L�����f�E�M�d�    Y_^[��]������������������������������������������U��Q�=,��u����=,��u���  �(j �E�Pj�MQ�,�R����u���  �f�E��]�����������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u�����     ��X��� 	   ����b  �} |�E;\�s	�E�   ��E�    �M��M܃}� u#h`hpjj jTh��j�.������u̃}� u9�j���     �xX��� 	   j jTh��h�h`��P���������  �E���M������P��D
��t	�E�   ��E�    �M؉Mԃ}� u#h�`hpjj jUh��j�������u̃}� u9�����     ��W��� 	   j jUh��h�h�`�(P��������5  �}���w	�E�   ��E�    �EЉẼ}� u#h$�hpjj jVh��j�	������u̃}� u9�E���     �SW���    j jVh��h�h$��O��������   �UR��[�����E�    �E���M������P��D
��t�MQ�UR�EP�0�����E��D��V��� 	   ����     �E�����3�u#h(ahpjj jah��j�:������u��E������   ��EP������ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   V�E�    �E������E��p����}�u�d���     �rU��� 	   �����  �} |�M;\�s	�E�   ��E�    �U��U��}� u&h`hpjj h�   h��j�������u̃}� u<�����     ��T��� 	   j h�   h��hL�h`�FM��������[  �M���U������P��L��t	�E�   ��E�    �U��U��}� u&h�`hpjj h�   h��j�������u̃}� u<�I���     �WT��� 	   j h�   h��hL�h�`�L��������  �}���w	�E�   ��E�    �M��M��}� u&h$�hpjj h�   h��j�������u̃}� u<����     ��S���    j h�   h��hL�h$��L��������*  �E�    �} t �E���M������P��D
��t3���  �} tǅt���   �
ǅt���    ��t����M��}� u&hl�hpjj h�   h��j�������u̃}� u<�����     �S���    j h�   h��hL�hl��NK��������c  �E���M������P��D
$�����E�M�M��}�t�}��&  �  �U��u	�E�   ��E�    �E��E��}� u&h`dhpjj h�   h��j��������u̃}� u<�-���     �;R���    j h�   h��hL�h`d�J��������  �U���s	�E�   ��E��E��M��Mh�   h��j�UR�~�����E�}� u��Q���    ����    ����;  jj j �EP�o2�����M���u������P��D1(�T1,�   �U��u	�E�   ��E�    �E��E��}� u&h`dhpjj h�   h��j��
������u̃}� u<����     �Q���    j h�   h��hL�h`d�eI��������z  �U����U�E�E�M�MԋU���E������P��T��H��  �E���M������P��D
��
��  �} ��  �M���U������P��MԊT��Eԃ��EԋM���M�U���U�E���M������P��D

�E���?  �M���U������P�¹   k� �D%��
�  �} �  �M���U�����P��   k� �EԊL
%��Uԃ��UԋE���E�M���M�U���E�����P��   k� �D%
�E����   �M���U������P�¹   �� �T%��
tk�} te�E���M�����P��   �� �EԊL%��Uԃ��UԋE���E�M���M�U���E�����P��   �� �D%
�UR�SH������tL�E���M������P��D
%�   t*��l���Q�U���E������P��R���E��}� tk�E��ubj �M�Q�U��R�E�P�M���U������P��Q�P��u!���E؋U�R������E������
  �E����E��   j �M�Q�UR�E�P�M���U������P��Q����t�}� |�U�;Uv^���E؃}�u#��M��� 	   ����M؉�E������
  �,�}�mu�E�    ��	  ��U�R�������E�������	  �E�E܉E�M���U������P��L��   ��	  �U���  �}� tE�E����
u:�U���E������P��T���E���M������P��T�8�M���U������P��L����U���E������P��L�E�E��M��M��U�U�9U��?  �E������   �U���E������P��T��@u:�E���M������P��D
���M���U������P��D��U��E���
�U����U��E����E��  �  �M����t!�E��M����E����E��M����M��  �U�E�L�9M�sG�U��B��
u�M����M��U��
�E����E���M��U����M����M��U����U��)  �E����E��E�    j �M�Qj�U�R�E���M������P��
P����u	���E؃}� u�}� u�M���U����U���   �E���M������P��D
��HtH�M��
u�U��
�E����E��,�M���U����U��E���M������P��E�D
�X�M�;M�u�U��
u�E�� 
�M����M��6jj�j��UR�]+������x�����|����E��
t�M���U����U������E�+E�E��M���#  �}� �  �U����U��E����   u�U����U��e  �E�   �E����X���u"�}��E�;E�r�M����M��UЃ��U��͋E����X��U��}� u��I��� *   �E������  �E���;E�u�M�MЉM���   �U���E������P��T��H��   �E���M������P��E�� �D
�M����M��}�|0�U���E�����P��   k� �M��	�L%�U����U��}�u0�E���M�����P��   �� �E�� �D%�M����M��U�+UЉU��"j�E��ؙRP�EP�)������x�����|����M�+M�M싕p�����R�EP�M�Q�U�Rj h��  ��E�}� u��P�� �����E�������  �E�+E�9E�t	�E�   ��E�    �M���U������P��M��L0�U���U��  �}� �  �E�E��M��M�E�+����U�B9E���   �M����uB�E���M������P��D
���M���U������P��D�   �   �U����t �M��U�f�f��M����M��U���U��]�E�+����M�TA�9U�sI�E��H��
u�U���U��
   �M�f��U����U���E��M�f�f��E����E��M���M������U�+U�����U��l  �}� tE�E����
u:�U���E������P��T���E���M������P��T�8�M���U������P��L����U���E������P��L�E�E��M��M�U�U�9U���  �E������   �U���E������P��T��@u:�E���M������P��D
���M���U������P��D��U��E�f�f�
�U����U��E���E��9  �/  �M����t#�E��M�f�f��E����E��M���M��  �U�E�L�9M�sN�U��B��
u�M���M��
   �E�f��M����M���U��E�f�f�
�U����U��E���E��  �M���M��E�    j �U�Rj�E�P�M���U������P��Q����u	���E؃}� u�}� u�   �E�f��M����M��6  �U���E������P��T��H��   �Ẽ�
u�
   �U�f�
�E����E��   �M̉Mĺ   �E�f��M����M��U���E������P��UĊ�T�Eă��EċM���U�����P��   k� �EĊ �D
%�M���U�����P��   �� �D%
�b�M�;M�u�Ũ�
u�
   �M�f��U����U��;jj�j��EP�$������x�����|����M̃�
t�   �E�f��M����M��,����U�+U�U�E�;Et�M�Q�]B�����}��u�U�U���EȉE��E�^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EP�MQ�UR�EP�.����]��������������������U��EPj �MQh�l�T	����]���������������������U���0�E�    3��EԉE؉E܉E��E�E�E�MЉM��} t	�E�   ��E�    �U��U�}� u&h��hpjj h�  hпj��������u̃}� u.��=���    j h�  hпhT�h���G6��������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]��������������������������������������������������������������������U��EP�MQ�URh�l������]�������������������U��EPj �MQh�2������]���������������������U��EP�MQ�URh�2�����]�������������������U��EPj �MQ�UR�����]����������������������U���H�E�    3��E��E��EĉEȉẺEЉEԍM��M��} t	�E�   ��E�    �U��U�}� u&h��hpjj h�   hпj��������u̃}� u1�<���    j h�   hпh4�h���W4��������k  �} t	�E�   ��E�    �M��M�}� u&hX�hpjj h�   hпj�8�������u̃}� u1�;���    j h�   hпh4�hX���3���������   �E��@B   �M��U�Q�E��M��U��B����EP�MQ�UR�E�P��;�����E��} u�E��   �M��Q���U�E��M�H�}� |"�U���  3Ɂ��   �M܋U�����M����U�Rj �3�����E܋E��H���M�U��E�B�}� |!�M��� 3�%�   �E؋M�����E����M�Qj �g3�����E؋E���]�����������������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP�MQ������]��������������U���0�E������E�    �} t	�E�   ��E�    �E�E��}� u&h�hpjj h9  hпj���������u̃}� u1�R9���    j h9  hпh,�h��1��������9  �} u�} u�} u3��   �} t�} v	�E�   ��E�    �U�U�}� u&h��hpjj h?  hпj�_�������u̃}� u1�8���    j h?  hпh,�h����0��������  �M;M��   �w8����U��EP�MQ�UR�E��P�MQh/2�&�����E��}����   �}�t^�}���tU�U��;UsJ�E���M+�9h�s�h��U���E���M+ȉM�U���Rh�   �E�M�TAR�������7���8"u
��7���M�������  �c�7����U��EP�MQ�UR�EP�MQh/2��%�����E�3ҋE�Mf�TA��}��u"�}�u�s7���8"u
�i7���U������o  �}� ��   �   k� 3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E��M���Qh�   �U��R������}��u}3�t	�E�   ��E�    �M܉M؃}� u&h��hpjj hf  hпj�D�������u̃}� u1�6��� "   j hf  hпh,�h����.��������   ����{�}�t]�}���tT�E���;EsI�M����U+�9h�s
�h��E���M����U+щUԋE���Ph�   �M��U�DJP������}� }	�E�������M��MЋEЋ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EPj �MQ�UR�EPh�l�#�����E��}� }	�E�������M��M��E���]�����������������������������U����EP�MQ�UR�EP�MQh�l�"�����E��}� }	�E�������U��U��E���]���������������������������U���H�E�    3��E��E��EĉEȉẺEЉEԍM��M��} t	�E�   ��E�    �U�U��}� u&h��hpjj h�   hпj�W�������u̃}� u1�3���    j h�   hпh��h����+��������  �} t�} u	�E�    ��E�   �M�M�}� u&hP�hpjj h�   hпj���������u̃}� u1�'3���    j h�   hпh��hP��r+��������8  �E��@B   �M��U�Q�E��M��}���?v�U��B�����E���M��A�UR�EP�MQ�U�R�U���E��} u�E���   �}� ��   �E��H���M�U��E�B�}� |!�M��� 3�%�   �E��M�����E����M�Qj �1+�����E��}��tY�U��B���E܋M��U܉Q�}� |"�E��� 3ҁ��   �U؋E�����U��
��E�Pj ��*�����E؃}��t�E�� 3ɋU�Ef�LP��M��y }�����������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EPj �MQ�UR�EPh�2�J�����E��}� }	�E�������M��M��E���]�����������������������������U����EP�MQ�UR�EP�MQh�2�������E��}� }	�E�������U��U��E���]���������������������������U���$�E������} t	�E�   ��E�    �E��E�}� u&h�hpjj h  hпj��������u̃}� u1��/���    j h  hпh��h��D(���������  �} t�} v	�E�   ��E�    �U��U�}� u&h��hpjj h  hпj��������u̃}� u1�t/���    j h  hпh��h���'��������x  �MQ�UR�EP�MQ�URh/2�}�����E��}� }b�   k� 3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R�f�����}��uz3�t	�E�   ��E�    �M�M��}� u&h��hpjj h  hпj��������u̃}� u.�e.��� "   j h  hпh��h���&��������l�}� |c�}�t]�}���tT�E���;EsI�M����U+�9h�s
�h��E���M����U+щU܋E���Ph�   �M��U�DJP�}�����E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP������]������������������U����  ���3ŉE�ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    �EP��d��������ǅ����    �n,����P����} tǅH���   �
ǅH���    ��H�����L�����L��� u&h�hpjj h  hx�j��������u̃�L��� uI�,���    j h  hx�hT�h��N$����ǅ,���������d����~�����,����8  �} tǅ@���   �
ǅ@���    ��@�����8�����8��� u&h��hpjj h  hx�j��������u̃�8��� uI�Z+���    j h  hx�hT�h���#����ǅ(���������d����������(����  ǅ����    ǅ����    ǅ����    ǅ����    ǅt���    �Uf�f�������������� ����U���U�� ��� �  ������ �  �������� |%��������x�������������0����
ǅ0���    ��0���������������������������������������D�����D�����  ��D����$��Rǅ����   ������Q�UR������P�  ���J  ǅ����    ������������������������������������ǅ����    ǅ��������ǅ����    ��  �������������������� ������������wj���������R�$��R���������������E���������������4���������������#�������ʀ   ����������������������e  ��������*u:�UR�t����������������� }���������������������ى������k�����
�������LЉ������  ǅ����    ��  ��������*u'�EP������������������ }
ǅ���������k�����
�������DЉ������  ��������������������I������������.�1  ���������R�$��R�U���lu�M���M��������   �����������������������   �M���6u+�E�H��4u�U���U������ �  �������   �M���3u(�E�H��2u�U���U������%����������S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    ������#�������� ���������������   �������D  ��������������������A������������7��
  ��������\S�$� S��������0  u�������� ������ǅ����   �EP�������f�������������� ��   ���������   �   k� ������ǅT���   ��T���s������T���Ƅ���� ��d�����,��P��d�����,��� �HtQ������R������P��#������}
ǅ����   ��   k� f������f������������������ǅ����   �s	  �UR� ����������������� t�������x u#�p�������������R�,	�����������d������%   t/�������Q������������� �+���������ǅ����   �(ǅ����    �������Q���������������������  ��������0  u�������� �������������uǅ4���������������4�����4����������EP�#������������������� ��   ������ u�p�������������������ǅ����    ���������������������;�����}O���������tB��d�����*��P�������P��+������t������������������������������   ������ u�t�������ǅ����   ������������������������������������������ t���������t��������������뾋�����+��������������2  �UR���������\����������   3�tǅ`���   �
ǅ`���    ��`�����<�����<��� u&h�hpjj h�  hx�j��������u̃�<��� uI��"���    j h�  hx�hT�h��6����ǅ$���������d����f�����$���� 	  �g  �������� t��\���f������f����\����������ǅ����   �-  ǅ����   �������� f��������������@������������������ǅt���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Yh�  hp�j������]  P�X����������������� t ��������������������]  ��t����
ǅ�����   �E���E�M�Q��A�������������d����(��P������Q������R������P��t���Q������R�����P�   k���0�P��Ѓ���������   t6������ u-��d����'��P������R�   k�	��0�R��Ѓ���������gu;��������   u-��d����\'��P������R�   ����0�Q��Ѓ����������-u!��������   ��������������������������P��������������  ��������@������ǅ����
   �   ǅ����
   �   ǅ����   ǅ����   �
ǅ����'   ǅ����   ��������   t8�   k� �0   f��������������Q�   �� f������ǅ����   �)ǅ����   ��������   t������   �������������� �  t�UR������������������   ������%   t�MQ�������������������   �������� tE��������@t�MQ�s���������������������UR�W���������������������@��������@t�MQ�.��������������������UR������3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ������������������ }ǅ����   �%���������������������   ~
ǅ����   �����������u
ǅ����    �   i��  ������������������������������������������ �������������   �������RP������R������P�b�����0�������������RP������Q������R����������������������9~���������������������������������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0�������������������� �a  ��������@��   ��������   t!�   k� �-   f������ǅ����   �V��������t!�   k� �+   f������ǅ����   �*��������t�   k� �    f������ǅ����   ������+�����+�������|�����������u������Q�UR��|���Pj �  ����P���Q������R�EP������Q������R�  ����������t'��������u������R�EP��|���Qj0�;  �������� ��   ������ ��   ��������������������x�����x����������x�������x�������� ��   ��d����Y!��P��d����M!��� �HtQ������R������P�Q������X�����X��� ǅ���������2������Q�UR������P��  ���������X����������X����(��P���R������P�MQ������R������P�  �������� |'��������t������R�EP��|���Qj �  �������� tj������R�������ǅ����    ������������������d����A���������M�3��������]��ABgB�B^CmC�CE�B�B�B�B�B�B �I 6D�D�CEE ��IYEGL[F�IvE�K�HtLL+G�KL�O   	
����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E�H��@t�U�z u�E����U�
�4�EP�MQ�!�����Ё���  u�E� ������M����E�]�������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�U������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��~�U�    �E�E��M���M�}� ~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������뛋E�8 u�M�U���]����������������������������������������������U���<�} t�} v	�E�   ��E�    �E�E��}� u#h^hpjj jh��j���������u̃}� u0�=���    j jh��hp�h^�	�����   �o  �} ��   �U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U�E�Ph�   �M��Q�]������} t	�E�   ��E�    �U�U�}� u#h�^hpjj jh��j��������u̃}� u0�c���    j jh��hp�h�^������   �  �M�M��U�U��}� v�E����t�U����U��E����E��܃}� ��   �M� �}�tH�}���t?�}v9�U��9h�s
�h��E��	�M���M��U�Rh�   �E��P�T���������t3�t	�E�   ��E�    �E܉E؃}� u#hP�hpjj j h��j���������u̃}� u0�S���    j j h��hp�hP�������   �  �U��E��
�U���EċM����M��U���U�}� t�E����E�t�ȃ}� ��   �M� �}�tH�}���t?�}v9�U��9h�s
�h��E��	�M���MԋU�Rh�   �E��P�<������ _��t3�t	�E�   ��E�    �EЉẼ}� u#hP_hpjj j*h��j���������u̃}� u-�;��� "   j j*h��hp�hP_������"   �p�}�th�}���t_�U+U���;UsQ�E+E����M+�9h�s�h��U���E+E����M+ȉMȋU�Rh�   �E+E��M�TR�O�����3���]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���L�U�M�}� t	�E�   ��E�    �E��E܃}� u&h��hpjj h>  h��j���������u̃}� u3�:���    j h>  h��h��h��������   �  �}� v	�E�   ��E�    �U؉Uԃ}� u&h��hpjj h?  h��j�d�������u̃}� u3����    j h?  h��h��h��������   �  �M�� �}��tH�}����t?�}�v9�U��9h�s
�h��E��	�M���MЋU�Rh�   �E��P��������} t	�E�   ��E�   �M�;M�v	�E�   ��E�    �UȉUă}� u&h �hpjj hA  h��j�w�������u̃}� u3��
��� "   j hA  h��h��h �������"   �)  �}r�}$w	�E�   ��E�    �M��M��}� u&h��hpjj hB  h��j���������u̃}� u3�E
���    j hB  h��h��h��������   �  �E�    �E�E��} t+�M��-�U����U��E����E��M�ًU�� �ډM�U�E��E�M3�RQ�EP�MQ������E�U3�PR�MQ�UR�@����E�U�}�	v�E��W�M���U����U���E��0�M���U����U��E����E��} w�} v�M�;M�r��U�;U���   �   k� �U��
 �E�;E�s	�E�   ��E�    �M��M��}� u&h��hpjj hf  h��j��������u̃}� u0����� "   j hf  h��h��h���0�����"   �E�E��  �M����M��U���E��M��U���M�U���E����E��M���M�U�;U�r�3���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�}�����]��������������������������U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP��   �E��j �MQ�UR�EP�MQ��   �E��E���]�����������������������������U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ�w   ��]��������������������U��j �EP�MQ�UR�U�M����]�������������������U��j �EP�MQ�UR�EP�   ]���������������������U���D�} t	�E�   ��E�    �E�E�}� u#h��hpjj jfh��j�.�������u̃}� u0����    j jfh��h��h����������   �Y  �} v	�E�   ��E�    �U��U܃}� u#h��hpjj jgh��j賾������u̃}� u0����    j jgh��h��h���V������   ��  �M� �}�tH�}���t?�}v9�U��9h�s
�h��E��	�M���M؋U�Rh�   �E��P�3������} t	�E�   ��E�   �M;M�v	�E�   ��E�    �UЉŨ}� u#h �hpjj jih��j�̽������u̃}� u0�!��� "   j jih��h��h ��o������"   ��  �}r�}$w	�E�   ��E�    �MȉMă}� u#h��hpjj jjh��j�K�������u̃}� u0����    j jjh��h��h����������   �v  �E�    �E�E��} t �M��-�U����U��E���E�M�ىM�U��U��E3��u�U�E3��u�E�}�	v�E��W�M���U����U���E��0�M���U����U��E���E�} v�M�;Mr��U�;U��   �   k� �U�
 �E�;Es	�E�   ��E�    �M��M��}� u&h��hpjj h�   h��j��������u̃}� u0�o��� "   j h�   h��h��h���������"   �E�E��  �M����M��U���E��M��U����M��U���E����E��M����M��U�;U�r�3���]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���L�U�M�}� t	�E�   ��E�    �E��E܃}� u&h��hpjj h>  h��j�E�������u̃}� u3� ���    j h>  h��h�h����������   �  �}� v	�E�   ��E�    �U؉Uԃ}� u&h��hpjj h?  h��j�Ĺ������u̃}� u3� ���    j h?  h��h�h���d������   �,  3ɋU�f�
�}��tK�}����tB�}�v<�E��9h�s�h��M��	�U���UЋE���Ph�   �M��Q�<������} t	�E�   ��E�   �U�;U�v	�E�   ��E�    �EȉEă}� u&h �hpjj hA  h��j�Ҹ������u̃}� u3�'���� "   j hA  h��h�h ��r������"   �:  �}r�}$w	�E�   ��E�    �U��U��}� u&h��hpjj hB  h��j�K�������u̃}� u3�����    j hB  h��h�h����������   �  �E�    �M�M��} t0�-   �E�f��M����M��U����U��E�؋M�� �ىE�M�U��U�E3�QP�UR�EP�L����E�M3�RQ�EP�MQ�����E�U�}�	v�U��W�E�f��M����M���U��0�E�f��M����M��U����U��} w�} v�E�;E�r��M�;M���   �   k� 3ɋU�f��E�;E�s	�E�   ��E�    �M��M��}� u&h��hpjj hf  h��j��������u̃}� u0�7���� "   j hf  h��h�h���������"   �M3��M�f��U����U��E�f�f�M��U��E�f�f�
�U�f�E�f��M����M��U���U�E�;E�r�3���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�m�����]��������������������������U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP��   �E��j �MQ�UR�EP�MQ��   �E��E���]�����������������������������U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ�w   ��]��������������������U��j �EP�MQ�UR�U�M�t���]�������������������U��j �EP�MQ�UR�EP�   ]���������������������U���D�} t	�E�   ��E�    �E�E�}� u#h��hpjj jfh��j�~�������u̃}� u0������    j jfh��h�h���!������   �o  �} v	�E�   ��E�    �U��U܃}� u#h��hpjj jgh��j��������u̃}� u0�X����    j jgh��h�h���������   ��  3ɋUf�
�}�tK�}���tB�}v<�E��9h�s�h��M��	�U���U؋E���Ph�   �M��Q�~������} t	�E�   ��E�   �U;U�v	�E�   ��E�    �EЉẼ}� u#h �hpjj jih��j��������u̃}� u0�l���� "   j jih��h�h ��������"   �  �}r�}$w	�E�   ��E�    �UȉUă}� u#h��hpjj jjh��j薱������u̃}� u0������    j jjh��h�h���9������   �  �E�    �M�M��} t%�-   �E�f��M����M��U���U�E�؉E�M��M��E3��u�U�E3��u�E�}�	v�U��W�E�f��M����M���U��0�E�f��M����M��U���U�} v�E�;Er��M�;M��   �   k� 3ɋUf��E�;Es	�E�   ��E�    �M��M��}� u&h��hpjj h�   h��j�\�������u̃}� u0����� "   j h�   h��h�h����������"   �M3��M�f��U����U��E�f�f�M��U��E�f�f�
�U�f�E�f��M����M��U����U��E�;E�r�3���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��} u�  �E�H;4�tj�U�BP�<������M�Q;8�tj�E�HQ�������U�B;<�tj�M�QR��������E�H;@�tj�U�BP�߼�����M�Q;D�tj�E�HQ��������U�B ;H�tj�M�Q R衼�����E�H$;L�tj�U�B$P肼�����M�Q8;`�tj�E�H8Q�c������U�B<;d�tj�M�Q<R�D������E�H@;h�tj�U�B@P�%������M�QD;l�tj�E�HDQ�������U�BH;p�tj�M�QHR�������E�HL;t�tj�U�BLP�Ȼ����]��������������������������������������������������������������������������������������������������������������U���VW�E�    �E�E��E�    �   k��E���    u�   ���U��
�    �n  jSh4�jjPj��������E��}� u
�   �  jYh4�jj�<������E�}� uj�E�P轺�����   ��  �M��    �   k��M���    �o  jeh4�jj�������E��}� u&j�U�R�g�����j�E�P�Y������   �u  �M��    �   k��M���   �U��E�    �E���Pj�M�Qj�U�R�������E��E��E���Pj�M�Qj�U�R������E��E��E���Pj�M�Qj�U�R������E��E��E���Pj�M�Qj�U�R�b�����E��E��E���Pj�M�Qj�U�R�A�����E��E��E��� PjP�M�Qj�U�R� �����E��E��E���$PjQ�M�Qj�U�R�������E��E��E���(Pj�M�Qj �U�R�������E��E��E���)Pj�M�Qj �U�R������E��E��E���*PjT�M�Qj �U�R������E��E��E���+PjU�M�Qj �U�R�{�����E��E��E���,PjV�M�Qj �U�R�Z�����E��E��E���-PjW�M�Qj �U�R�9�����E��E��E���.PjR�M�Qj �U�R������E��E��E���/PjS�M�Qj �U�R�������E��E��E���8Pj�M�Qj�U�R�������E��E��E���<Pj�M�Qj�U�R������E��E��E���@Pj�M�Qj�U�R������E��E��E���DPj�M�Qj�U�R�s�����E��E��E���HPjP�M�Qj�U�R�R�����E��E��E���LPjQ�M�Qj�U�R�1�����E��E�t@�E�P耼����j�M�Q�Y�����j�U�R�K�����j�E�P�=������   �Y  �M��QR�  ����   �(��}��E���   �U����M���   �E��J�H�U���   �M��P�Q�E���   �U��A0�B0�M���   �E��J4�H4�U��   �}� t	�E��    ��E�    �E�    �E�(��M���    tE�U���   �����Iu2�U���    w&hd�hpjj h�   h��j蛧������u̋M�yx t5�U�Bx�����Iu%j�U���   P������j�M�QxR��������E�M����   �U�E�Bx�M�U����   3�_^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]������������������������������������U��} u�   �E�;(�tj�U�P螳�����M�Q;,�tj�E�HQ�������U�B;0�tj�M�QR�`������E�H0;X�tj�U�B0P�A������M�Q4;\�tj�E�H4Q�"�����]��������������������������������������������������������U���VW�E�    �E�    �E�E��E�    �   ���U��
�    u�   k��U��
�    �1  jeh�jjPj�[������E��}� u
�   ��  �E�   ���   �}��jqh�jj貟�����E��}� uj�M�Q�3������   �}  �U��    �   ���M���    �E  j}h�jj�\������E�}� u&j�U�R�ݱ����j�E�P�ϱ�����   �  �M��    �   ���E���   �M�U�Rj�E�Pj�M�Q�E�����E��E��U���Rj�E�Pj�M�Q�$�����E��E��U���Rj�E�Pj�M�Q������E��E��U���0Rj�E�Pj�M�Q�������E��E��U���4Rj�E�Pj�M�Q�������E��E�t0�U�R�޵����j�E�P������j�M�Q�۰��������'  �U��BP��  ���A�E�    �M��(���E��,��H�U��0��B�M��X��Q0�E��\��H4�U��   �}� t	�E��    ��E�    �E�    �E�(��M�y| t?�U�B|�����Iu/�U�z| w&h@�hpjj h�   h��j�j�������u̋M�yx t5�U�Bx�����Iu%j�U�BxP������j�M���   R�̯�����E�M�H|�U�E��Bx�M�U����   3�_^��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]������������������������������������U��} u�	  j�   �� �M�R������j�   ���M�R������j�   k��U�
P�ѭ����j�   ���U�
P踭����j�   k��E�Q蟭����j�   k��M�R膭����j�   k� �U�
P�m�����j�   �� �U�D
P�S�����j�   ��U�D
P�:�����j�   k��E�LQ� �����j�   ���E�LQ������j�   k��M�TR������j�   k��U�D
P�Ҭ����j�   k� �E�LQ踬����j�   k� �M�T8R螬����j�   �� �M�T8R脬����j�   ���M�T8R�k�����j�   k��U�D
8P�Q�����j�   ���U�D
8P�7�����j�   k��E�L8Q������j�   k��M�T8R������j�   k��U�D
8P������j�   ���U�D
8P�ϫ����j�   k�	�E�L8Q赫����j�   k�
�M�T8R蛫����j�   k��U�D
8P聫����j�   k� �E�LhQ�g�����j�   �� �E�LhQ�M�����j�   ��E�LhQ�4�����j�   k��M�ThR������j�   ���M�ThR� �����j�   k��U�D
hP������j�   k��E�LhQ�̪����j�   k��M�ThR貪����j�   ���M�ThR蘪����j�   k�	�U�D
hP�~�����j�   k�
�E�LhQ�d�����j�   k��M�ThR�J�����j�   k� �U��
�   P�-�����j�   �� �U��
�   P������j�M���   R�������j�E���   Q������j�U���   P�ԩ����j�   �� �U��
�   P跩����j�   ��U��
�   P蛩����j�   k��E���   Q�~�����j�   ���E���   Q�a�����j�   k��M���   R�D�����j�   k��U��
�   P�'�����j�   k� �E���   Q�
�����j�   �� �E���   Q������j�   ��E���   Q�Ѩ����j�   k��M���   R质����j�   ���M���   R藨����j�   k��U��
�   P�z�����j�   k��E���   Q�]�����j�   k� �M���   R�@�����j�   k� �U��
�   P�#�����j�   �� �U��
�   P������j�   ��U��
�   P������j�   k��E���   Q�ͧ����j�   ���E���   Q谧����j�   k��M���   R蓧����j�   k��U��
�   P�v�����j�   k��E���   Q�Y�����j�   ���E���   Q�<�����j�   k�	�M���   R������j�   k�
�U��
�   P������j�   k��E���   Q������j�   k� �M��  R�Ȧ����j�   �� �M��  R諦����j�   ���M��  R菦����j�   k��U��
  P�r�����j�   ���U��
  P�U�����j�   k��E��  Q�8�����j�   k��M��  R������j�   k��U��
  P�������j�   ���U��
  P������j�   k�	�E��  Q�ĥ����j�   k�
�M��  R觥����j�   k��U��
  P芥����j�   k� �E��L  Q�m�����j�   �� �E��L  Q�P�����j�U��T  P�<�����j�M��X  R�(�����j�E��\  Q������j�U��`  P� �����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�   k��U��
�    trj@h��jhd  j�P������E��}� u
�   �   �EP�M�Q��   ����t$�U�R�x�����j�E�P�7������   �   �M�ǁ�      ��E����U���   ��tN�E���   ���   �����Ju5�E���   ���    #h �hpjj jPhx�j��������u̋E�M����   3���]��������������������������������������������������������������������������������U����E�    �   k��U��
�   �E��   k��E���   �M�} u����  �U�R�������M��`  �U�U��E�    �   �� EPj1�M�Qj�U�R舽����E��E��   ��EPj2�M�Qj�U�R�c�����E��E��   k�MQj3�U�Rj�E�P�=�����E��E��   ��MQj4�U�Rj�E�P������E��E��   k�URj5�E�Pj�M�Q������E��E��   k�EPj6�M�Qj�U�R�˼����E��E��   k� MQj7�U�Rj�E�P襼����E��E��   �� �U�D
Pj*�M�Qj�U�R�{�����E��E��   ���M�TRj+�E�Pj�M�Q�R�����E��E��   k��M�TRj,�E�Pj�M�Q�(�����E��E��   ���E�LQj-�U�Rj�E�P�������E��E��   k��E�LQj.�U�Rj�E�P�Ի����E��E��   k��E�LQj/�U�Rj�E�P誻����E��E��   k� �E�LQj0�U�Rj�E�P耻����E��E��   k� �E�L8QjD�U�Rj�E�P�V�����E��E��   �� �U�D
8PjE�M�Qj�U�R�,�����E��E��   ���M�T8RjF�E�Pj�M�Q������E��E��   k��M�T8RjG�E�Pj�M�Q�ٺ����E��E��   ���E�L8QjH�U�Rj�E�P诺����E��E��   k��E�L8QjI�U�Rj�E�P腺����E��E��   k��E�L8QjJ�U�Rj�E�P�[�����E��E��   k��E�L8QjK�U�Rj�E�P�1�����E��E��   ���U�D
8PjL�M�Qj�U�R������E��E��   k�	�U�D
8PjM�M�Qj�U�R�ݹ����E��E��   k�
�U�D
8PjN�M�Qj�U�R賹����E��E��   k��U�D
8PjO�M�Qj�U�R艹����E��E��   k� �U�D
hPj8�M�Qj�U�R�_�����E��E��   �� �M�ThRj9�E�Pj�M�Q�5�����E��E��   ��E�LhQj:�U�Rj�E�P������E��E��   k��E�LhQj;�U�Rj�E�P������E��E��   ���U�D
hPj<�M�Qj�U�R踸����E��E��   k��U�D
hPj=�M�Qj�U�R莸����E��E��   k��U�D
hPj>�M�Qj�U�R�d�����E��E��   k��U�D
hPj?�M�Qj�U�R�:�����E��E��   ���M�ThRj@�E�Pj�M�Q������E��E��   k�	�M�ThRjA�E�Pj�M�Q������E��E��   k�
�M�ThRjB�E�Pj�M�Q輷����E��E��   k��M�ThRjC�E�Pj�M�Q蒷����E��E��   k� �M���   Rj(�E�Pj�M�Q�e�����E��E��   �� �E���   Qj)�U�Rj�E�P�8�����E��E��M���   Qj�U�Rj�E�P������E��E��M���   Qj �U�Rj�E�P������E��E��M���   Qh  �U�Rj�E�P�ɶ����E��E��M���   Qh	  �U�Rj �E�P袶����E��E��   �� �U��
�   Pj1�M�Qj�U�R�u�����E��E��   ���M���   Rj2�E�Pj�M�Q�I�����E��E��   k��M���   Rj3�E�Pj�M�Q������E��E��   ���E���   Qj4�U�Rj�E�P������E��E��   k��E���   Qj5�U�Rj�E�P�µ����E��E��   k��E���   Qj6�U�Rj�E�P蕵����E��E��   k� �E���   Qj7�U�Rj�E�P�h�����E��E��   �� �U��
�   Pj*�M�Qj�U�R�;�����E��E��   ���M���   Rj+�E�Pj�M�Q������E��E��   k��M���   Rj,�E�Pj�M�Q������E��E��   ���E���   Qj-�U�Rj�E�P赴����E��E��   k��E���   Qj.�U�Rj�E�P舴����E��E��   k��E���   Qj/�U�Rj�E�P�[�����E��E��   k� �E���   Qj0�U�Rj�E�P�.�����E��E��   k� �E���   QjD�U�Rj�E�P������E��E��   �� �U��
�   PjE�M�Qj�U�R�Գ����E��E��   ���M���   RjF�E�Pj�M�Q訳����E��E��   k��M���   RjG�E�Pj�M�Q�{�����E��E��   ���E���   QjH�U�Rj�E�P�N�����E��E��   k��E���   QjI�U�Rj�E�P�!�����E��E��   k��E���   QjJ�U�Rj�E�P�������E��E��   k��E���   QjK�U�Rj�E�P�ǲ����E��E��   ���U��
�   PjL�M�Qj�U�R蚲����E��E��   k�	�U��
�   PjM�M�Qj�U�R�m�����E��E��   k�
�U��
�   PjN�M�Qj�U�R�@�����E��E��   k��U��
�   PjO�M�Qj�U�R������E��E��   k� �U��
  Pj8�M�Qj�U�R������E��E��   �� �M��  Rj9�E�Pj�M�Q蹱����E��E��   ��E��  Qj:�U�Rj�E�P荱����E��E��   k��E��  Qj;�U�Rj�E�P�`�����E��E��   ���U��
  Pj<�M�Qj�U�R�3�����E��E��   k��U��
  Pj=�M�Qj�U�R������E��E��   k��U��
  Pj>�M�Qj�U�R�ٰ����E��E��   k��U��
  Pj?�M�Qj�U�R謰����E��E��   ���M��  Rj@�E�Pj�M�Q������E��E��   k�	�M��  RjA�E�Pj�M�Q�R�����E��E��   k�
�M��  RjB�E�Pj�M�Q�%�����E��E��   k��M��  RjC�E�Pj�M�Q�������E��E��   k� �M��L  Rj(�E�Pj�M�Q�˯����E��E��   �� �E��L  Qj)�U�Rj�E�P螯����E��E��M��T  Qj�U�Rj�E�P�z�����E��E��M��X  Qj �U�Rj�E�P�V�����E��E��M��\  Qh  �U�Rj�E�P�/�����E��E��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��SVWUj j h���u�����]_^[��]ËL$�A   �   t2�D$�H�3�荞��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h��d�5    ���3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y��u�Q�R9Qu�   �SQ����SQ����L$�K�C�kUQPXY]Y[� ��������������������������������������������������������������������������������������������U��Q�M��E��     �E���]����������U����M��E��H�� ����U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M�9 ��  �U������  �E�    �U��E���M����E��M�����  �M���M;���   �U����_��   �U����$��   �U����<��   �U����>��   �U����-tw�U����a|�U����z~]�U����A|�U����Z~C�U����0|�U����9~)�U�����   |�U�����   ~	��v����t�U����U���E��H�� ������U��J�   ������E�P�M�Q�M�������U����tG�U���M��U�U�E����U�
�E�;E�t�M��Q�� ������E��P�M��    � �M�赢����u�U��B% ������M��A��U��B% ������M��A��U��B% ������M��A�E���]� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M��E��M���I�H�E���]� ����������������U��Q�M��E��H�� ����U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M�衱���E���]� ���������������������������������������������������������������U����M��} tpj h`�j�l������E��}� t�EP�M������E���E�    �M��U��E��8 t	�E�    ��E�   �M����   �U��B% �����M��A��U��B% ����M��A�U��    �E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E���]� ������������������������������������������������������������������������������U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} t%�MQ�m�  ���E��}� v�U�R�EP�M�������E���]� ������������������������������������������������������������������������U����M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�}t�}t	�E�    ��E�E��M����   �U��B% �����M��A�U��    �}u.�EP��������M���U��: u�E��H�� ������U��J�E���]� ��������������������������������������������������������������������������U��Q�M��E��     �M��Q�� ����E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�E���]��������������������������������������������������������U���(���3ŉE��M��E��E؋M��Q�� ����E��P�M��    �U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%����M��A�U�� �E� �} |�} s�E��E�؋M�� �ىE�M�U؃��U�j j
�EP�MQ�;�����0�� �U؈j j
�EP�MQ耋���E�U�UUu��E߅�t�M؃��M؋U��-�E؍M�+��   +�R�E�P�M�������E��M�3��������]� �����������������������������������������������������������������������������������������������������������U���$���3ŉE��M��E��E܋M��Q�� ����E��P�M��    �U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%����M��A�U�� �E܃��E�j j
�MQ�UR脋����0�� �M܈j j
�UR�EP�ɉ���E�U�MMu��U܍E�+й   +�Q�U�R�M��W����E��M�3��^�����]� �������������������������������������������������������������������������������������������U��Q�M��E�� ��E���]����������U����M��M��O����E�� l��M��U�Q�E��xu	�E�   ��E�    �M��U��Q�E���]� ����������������������������������U��Q�M��E�� �����E���]����������U��Q�M��M��X����M���,�M����E�H��H��D��} t�U�P��E�L���L�    �P�    �M���,�<��U��8��E�T��M�\��X� �E���]� �����������������������������������������������U��Q�M��M������E�� 0��M��U�Q�E���]� ����������������������U����M��M�迃���E�� X��} t#�M�,�����t�M������u	�E�    ��M�M��U��E��B�E���]� �������������������������������������U��Q�M��M��A����E�� ���M��U�Q�E��M�H�U��B�����E���]� �������������������U����M��M������E�� D��} t\�} tVj h`��MQ�c{�����E��U��E��B�M��U�Q�E��x t�MQ�UR�E��HQ��  ���
�U��B    ��E��@    �M��A    �E���]� ���������������������������������������U��EP�MQ�`��x���]����������U��Q�M��E��M���I�H�E���]� ����������������U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M�葤���E���]� ���������������������������������������������������������������U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} tXj h`�j�x�����E��}� t�MQ�M��)����E���E�    �U��E��M��9 u�U��B% ������M��A��U��B% ������M��A�E���]� ���������������������������������������������������������������������������������U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�MQ�e�  ��P�UR�M�������E���]� ������������������������������������������������������������U��Q�M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E%�   �M��Q�� ���ЋE��P�}u0�MQ�1������U���E��8 u�M��Q�� ������E��P�	�M��    �E���]� ���������������������������������������������������������������������U��Q�M��} |�}	~j�M蹢���E�;�9�E��8�t
�M��U;~j�M薢���E���E�M��T�R�M�dt���E��]� �����������������������������U���H�M��M��x����M��p����=H� �E  �H����?uQ�   �� �H����@u;�D����D��E�P��l����PhL��M�Q�^w����P�M��%c����   �H����?ut�   �� �H��
��$u]j �M�Q�[z����P�M���b���M��L�����t�z����u.�D����t!�H��D��U�R�Wl����P�M��b���e�   k� �H��
��?u9�   �� �H��
��?u"�   ��H��
��@uj�M�������M�Q��k����P�M��9b���M�衍����u	3��  �@�M�苍����t��y����u�D����t�H�Q�M��9�����U�R�M���a���=L� u1�M��V������P�jh`��P�P�=s�����E�M�L��=L� ��   �P�R�L�P�M��^����L��M��U��U��E����tY�U���� u0�M����M��U�� �E����E��M���� u�E����E�����M��U����M����M��U����U�띋E��M����L���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EP�MQ�UR�M�趡����萉���E��]������������������������U����EP�MQ�UR�M��������Q����E��]�������������������������U����EP�MQ�UR�M��l����������E��]�������������������������U����M��E�P�M��p���MQ�M�菱���U�R�M�p���E��]� ��������������������������U����M��E�P�M���o���MQ�M������U�R�M�o���E��]� �������������������������U����M��E�P�M��yo���MQ�M��k����U�R�M�ao���E��]� ��������������������������U����M��E�P�M��)o���MQ�M�������U�R�M�o���E��]� ��������������������������U����M��E�P�M���n���MQ�M��`����U�R�M��n���E��]� ��������������������������U��Q�M��M��k����tG�M�k����t�M�M���P�M������(�M��k����t�EP�M��]����M�R�M���r���E���]� �����������������������������U����M��M��j����tb�E��tZ�M��k����t�MQ�M���t���?j h`�j��n�����E��}� t�UR�M��J����E���E�    �E�P�M��4r���E���]� ��������������������������������U����M��M���i������   �} ��   �M��tj����t�EP�M��zc���j�M������t�M������u@j h`�j�n�����E��}� t�MQ�M��}����E���E�    �U�R�M��wq����M趇��P�M��j����E���]� ������������������������������������������������U����M��M��i����tu�} to�E���te�M��i����t�UR�M������Kj h`�j�<m�����E��}� t�EP�N�  ��P�MQ�M��\����E���E�    �U�R�M��p���E���]� ���������������������������������������������U��Q�M��M��_h����tC�M���h����u�}t�}u�EP�M��̂����} u��MQ�v����P�M��p���E���]� ���������������������������������U����M��M��]����uj�M�bh����u^j h`�j�l�����E��}� t�EP�M��k���E���E�    �M�M�}� t �U�����E��M��U���E��M��U�T��E���]� ����������������������������������������U����M��M��s�����t3�M� g����u'�M�Z����E��E�%�   �M��Q�� ���ЋE��P�E���]� ������������������������������U��Q�M��E��M��U��E�B�M��A    �U��B    �E��@    ��]� ��������������������U��Q�M��E��x t7�M��U��B�A�M��y t"�U��B�M���Q�E��HQ�U��B�Ѓ��ɋ�]����������������������U���l�����t�E�������M������]������������������������U����M��} t_j h`�j�j�����E��}� t�EP�M��R�M��h���E���E�    �E��M��U��: u�E��H�� ������U��J��E��H�� ������U��J��]� ���������������������������������������U���  �M��؆�������E��M��\���������}���  uj�M�|����E�8  �B�}���  u�EPj�MQ�E������E�  ��}���  u�UR�M� h���E��  �E�% �  �{  �M��� �  t5�U���   ��   uǅt���   �
ǅt���    ��t����������-�M��� `  uǅ����   �
ǅ����    ������������������ t�E�%   �E���M���   �M��}� tL�U��� �  t0�E�%   =   uǅ����   �
ǅ����    �������M���E�    �}� ��  �U��� �  t3�E�%   =   uǅ����   �
ǅ����    �������������$�U��� `  u	�E�   ��E�    �EЉ����������� t�M���   �M���U���   �Uȃ}� ��   �E�% �  t2�M���   ��   uǅ����   �
ǅ����    �������U���E�    �}� ��  �E�% �  t2�M���   ��   uǅ����   �
ǅ����    �������U���E�    �}� �q  �E�% @  tV�X����t5蚁����t,��p���Q�^����Pj ��`���R�`�����P�M�� U���������P��]����P�M��o���M��� �  t5�U���   ��   uǅ����   �
ǅ����    �������������$�M��� `  u	�E�   ��E�    �U������������� t�E�%   �E���M���   �M��}� �O  �U��� �  t0�E�%   =   uǅ����   �
ǅ����    �������M���E�    �}� �  ������R�e����P������Pj{�����Q�M��{�����Y}��P�M�����������R�������k����u4h����p���P������Qj,������R���������d���P�M��¥��h���M�����������P��y������V����tU��y����tL�)k����uC�M�Q��`���Rj ��P���P������Qj ��P���R�z��������{�����|��P�M��,S���-
  �������������������������������������������������Ձ���E�% �  t5�M���   ��   uǅ����   �
ǅ����    �������������#�E�% `  u	�E�   ��E�    �M������������� t�U���   �U���E�%   �E��}� ��  �M��� �  t5�U���   ��   uǅ����   �
ǅ����    �������������$�M��� `  u	�E�   ��E�    �U������������� te�E�%   =   uV������Q�.q����P��������Q����@���R�q����P�������Q���� ���P��p����P�������Q���   �M��� �  t,�U���   ��   u	�E�   ��E�    �E���x����-�M��� `  uǅ����   �
ǅ����    ��������x�����x��� t*�E�%   =   u��0���Q�\p����P��������P��������R�Ap����P��������P���E�% �  t5�M���   ��   uǅ����   �
ǅ����    ��������x����,�E�% `  uǅp���   �
ǅp���    ��p�����x�����x��� �  �U��� �  t3�E�%   =   uǅh���   �
ǅh���    ��h�����`����-�U��� `  uǅp���   �
ǅp���    ��p�����`�����`��� tS�M��� �  t5�U���   ��   uǅh���   �
ǅh���    ��h�����X����
ǅX���   ��X��� uA�
�����t�� ���Q�X�����P�������{O�����@���R�;�����P�������li���R����tO�u����t,�E�P�����Q������R�u�������x��P�M��"O����� ���P�u����P�M��i����� ���Q�eu����P�M���h���M�\����uA�M��\����u)�f����u �URj ������P������P�M��ˠ����MQ�M��N���E�    �������t}�������� tNj ������R��}����PhT�������P�b����P�M��s����f����t�M�Q�M��^���E�  �ej h`�j�_������`�����`��� t��`�����|����P����
ǅP���    ��P����U��E�P��0���Q�g}����P��������M���U��� �  t3�E�%   =   uǅX���   �
ǅX���    ��X�����P����-�U��� `  uǅH���   �
ǅH���    ��H�����P�����P��� t�M���   ��@�����U���   ��@�����@��� ��  �E�% �  t5�M���   ��   uǅH���   �
ǅH���    ��H�����@����,�E�% `  uǅ8���   �
ǅ8���    ��8�����@�����@��� ��   �U���   ��   ��   j,������P������Q������Rj,������P������Q������Rj,��x���P������Qh����h���R�`�������.t�����u����� t�����u�����t��P�M��C�����   �E�% �  t5�M���   ��   uǅ0���   �
ǅ0���    ��0�����(����,�E�% `  uǅ8���   �
ǅ8���    ��8�����(�����(��� tG�U���   ��   u6j,��X���P������Qh���H���R�_�������Ts��P�M�腝���h��M��Վ��h����8���P�����������P�M��V���j)��(���Q�����R�bc����Pj(�����P�G���������r��P�M������M��� �  t5�U���   ��   uǅ0���   �
ǅ0���    ��0�����(����-�M��� `  uǅ ���   �
ǅ ���    �� �����(�����(��� ��   �E�% �  t5�M���   ��   uǅ���   �
ǅ���    �����������,�E�% `  uǅ ���   �
ǅ ���    �� ������������� tQ�U��� �  t3�E�%   =   uǅ���   �
ǅ���    �����������
ǅ���   ����� u������R�M��Λ���U�����t������P�O[����P�M�譛���������Q�5[����P�M��c���V����t������R�}����P�M��r����������P�i}����P�M��Jc��������Q��y����P�M��2c���'n����t!�}� t�U�R�M��	I��������P�M���H����  �MQ�M������U��� �  u,�E�% |  = h  u�M�Q�UR�6\�����E�-  �  �E�% �  u.�M��� |  �� p  u�U�R�EP�L�����E��  ��  �M��� �  u]�U��� |  �� `  uLh���EP������Q�ZU����P������Rj{������P�M��p�����q������~���E�  �g  �M��� �  u.�U��� |  �� |  u�E�P�MQ�S�����E�T  �.  �U��� �  t3�E�%   =   uǅ���   �
ǅ���    �����������-�U��� `  uǅ ���   �
ǅ ���    �� ������������� t�M���   ��������U���   ������������ td�E�% �  t5�M���   ��   uǅ ���   �
ǅ ���    �� ����������
ǅ����    ������ th,��M��X����-  �E�% �  t5�M���   ��   uǅ����   �
ǅ����    �������������,�E�% `  uǅl���   �
ǅl���    ��l��������������� t�U���   ��,�����E�%   ��,�����,��� te�M��� �  t5�U���   ��   uǅ����   �
ǅ����    ��������d����
ǅd���    ��d��� thT��M��W����,  �M��� �  t5�U���   ��   uǅ����   �
ǅ����    �������������-�M��� `  uǅ���   �
ǅ���    ����������������� t�E�%   ��\�����M���   ��\�����\��� t`�U��� �  t3�E�%   =   uǅ����   �
ǅ����    ��������$����
ǅ$���    ��$��� th���M��V����.�U��� �  u#�E�% |  = x  u�M�Q�M�MU���E�!	  �U��� �  t3�E�%   =   uǅ����   �
ǅ����    �������������-�U��� `  uǅT���   �
ǅT���    ��T��������������� t�M���   ��������U���   ������������ ��   �E�% �  t5�M���   ��   uǅ����   �
ǅ����    ��������L����
ǅL���    ��L��� uR�E�% �  t5�M���   ��   uǅ����   �
ǅ����    ������������
ǅ���    ����� t#�E�PhT���x���Q�~W����P�M��EC����U�R��h���P�R����P�M��'C���M��� �  t5�U���   ��   uǅ����   �
ǅ����    �������������-�M��� `  uǅD���   �
ǅD���    ��D��������������� �#  �&`�����   �E�% �  t5�M���   ��   uǅ���   �
ǅ���    �������<����,�E�% `  uǅ����   �
ǅ����    ��������<�����<��� tr�U��� �  t3�E�%   =   uǅ����   �
ǅ����    ������������
ǅ���   ����� t!�U�Rh����X���P��U����P�M��A���M��� �  t�U���   ��   ��  �E�% �  t2�M���   ��   uǅ|���   �
ǅ|���    ��|����U��)�E�% `  uǅ4���   �
ǅ4���    ��4����M�}� t�U���   ��������E�%   ������������ �c  �M��� �  t)�U���   ��   u	�E�   ��E�    �E�E��!�M��� `  u	�E�   ��E�    �U�U܃}� t�E�%   =   ��   �M��� �  t)�U���   ��   u	�E�   ��E�    �EԉE��!�M��� `  u	�E�   ��E�    �ỦUă}� t�E�%   =   tj�M��� �  t)�U���   ��   u	�E�   ��E�    �E��E��!�M��� `  u	�E�   ��E�    �U��U��}� t0�E�%   =   u!�M�Qh����H���R��S����P�M��?���	������	  �E�% �  t)�M���   ��   u	�E�   ��E�    �U��U�� �E�% `  u	�E�   ��E�    �M��M��}� ��   �U��� �  t(�E�%�   ��@u	�E�   ��E�    �M���|����*�U���   ��   u	�E�   ��E�    �E���|�����|��� t&�M�Qh����8���R��R����P�M��>���   �E�% �  t5�M���   ��   uǅt���   �
ǅt���    ��t�����d����,�E�% `  uǅl���   �
ǅl���    ��l�����d�����d��� ��   �U��� �  t3�E�%�   =�   uǅ\���   �
ǅ\���    ��\�����L����3�U���   ��   uǅT���   �
ǅT���    ��T�����L�����L��� t&�M�Qh����(���R��Q����P�M��=���  �E�% �  t5�M���   ��   uǅD���   �
ǅD���    ��D�����4����,�E�% `  uǅ<���   �
ǅ<���    ��<�����4�����4��� ��   �U��� �  t.�E�%�   uǅ,���   �
ǅ,���    ��,���������-�U���   uǅ$���   �
ǅ$���    ��$������������� t!�M�Qh ������R��P����P�M��<���E�% �  t5�M���   ��   uǅ���   �
ǅ���    �����������,�E�% `  uǅ���   �
ǅ���    ��������������� t�U���   ��������E�%   ������������ t*�S����u!�M�Qh������R��O����P�M���;���E�%   t!�M�Qh�������R��O����P�M��;���E�P�M�'L���E��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M�jPh���M��%v�������]������������������U��Q�T�%�   u	�E�   ��E�    �E���]����������U��Q�T���u	�E�   ��E�    �E���]������������U��Q�T���u	�E�   ��E�    �E���]������������U��Q�T�% �  u	�E�   ��E�    �E���]����������U��Q�T�%   u	�E�   ��E�    �E���]����������U��Q�T���u	�E�   ��E�    �E���]������������U��Q�T���u	�E�   ��E�    �E���]������������U��Q�T�%   u	�E�   ��E�    �E���]����������U��T�%   ]������������������U��T�%   ]������������������U����M��E��8 tj�M��Z���  �} ��   �} ��   �M�M��}� t�}�t�u�U��B% ������M��A�   j h`�j�C�����E�}� t�U�P�M��v���E���E�    �M��U���E��8 u�M��Q�� ������E��P�[j h`�j�.C�����E�}� t�MQ�UR�M��Wg���E���E�    �E��M��U��: u�E��H�� ������U��J��E��H�� ������U��J��]� �������������������������������������������������������������������������������������������U��Q�T�%   u	�E�   ��E�    �E���]����������U��Q�T�%   u	�E�   ��E�    �E���]����������U��Q�T���`��`t	�E�   ��E�    �E���]�������������������������U��Q�T�%   u	�E�   ��E�    �E���]����������U��T�%    ]������������������U��Q�T���u	�E�   ��E�    �E���]������������U���,�E�   �M��^���M��[�����  �D����@��   �D����Z��   �}� t	�E�    �
j,�M��-Q���D������   �D����0�M�x3�}�	-�D����D��E�P�M�Q�8���1��P�M��-����k�D��U�M���]��P�E�P�bW�����D�+M��~�8��:1����u�U�R�8��k.���E�P�M��Հ���D�;M�u
j�M��cV���j�M���~���������U�R�M�?���E��]�������������������������������������������������������������������������������������������U��� �D���M��}�XtD�}�Zt�`�D����D��tV����t	�E�P��E���E�P�M��{���E��   �D����D�h���M��{���E��   �U�R�,S�����M��Y������   �D���M��}� t�}�@t`�}�Zt�v�U�R�M��=���E�   �D����D���U����t	�E����E���M�Q�U�R�M���c��P�M�=���E�>�D����D��M�Q�M�=���E� j�M�k���E���U�R�M�s=���E��]�����������������������������������������������������������������������������������������������U���   �D�����~  ��6���E��}� }�E�    �}� u>j]�U�Rj�E�Pj[�M��m�����L������S��P�MQ�@?�����E��  �   �M���Z���M�Df����th���M��\o���M��9����tZ�U��U��E����E��}� tE�D����t8j]��x���Pj �M�Q�h����Pj[�U�R��`�������hS��P�M��}��뚋M�.9����ua�M�e����t�E�P�M�Q�M�T��P�M��J+���:�U�R��h���Pj)�M�Q�URj(�E�P�\`������� S�����uT��P�M��+���M�Q�U�R�oS�����M��aL���E�P�M�;���E�   �   �M�8����uPj]�M�Qj�U�Rh ��E�P�MQj(�U�R��_�������Xa�����0K�����wR��P�EP�=�����E�<�:j]�M�Qj��p���Rj[��`�����k������J�����9R��P�EP�{=�����E��]������������������������������������������������������������������������������������������������������������������������������������������������U���j �X����P�M��w���D����tl�D���E��D����D��U��U��}�0t�}�2t�}�5t(�5h���M���l���&�E�P�y8����P�M��R{���j�M��g���E�(�
j�M��Fy��h(��M��l���M�Q�M�9���E��]������������������������������������������������������U���t�D�����k  �D���E��D����D��E� �E������M��fW���U��U�E��C�E�}��   �M�����$���h���M��]���?  h���M��]���-  h���M��m]���  h���M��[]���	  h���M��I]����  hD��M��7]��h���M��]k����  �E����E���  �D���U��E��E�D����D��U�U�}�Y�8  �E���\��$�(��E������(  h���M��\���  h���M��\���  h���M��\����   h��M��\����   h��M��s\����   h ��M��a\���   h,��M��O\���   h8��M��=\���   �D����D��E�P�+.����P�M���&���M��4����t�M�Q�M�N7���E�~  �R�UR�E�P��9����PhD��MQ�:�����E�R  �D����D�j�M��&N���hL��M��[���Qh���M��[���B�D����D��M�Q�-����P�M��%&���M���3����t�U�R�M�6���E��  �}����   �E��E��M���C�M��}���   �U������$����M�QhL��U�R��9����P�M��%���e�E�PhX��M�Q��9����P�M��%���E�U��U�E��E�E�}�w/�M������$����E�PhL��M�Q�9����P�M��K%���M��2����u�URj �E�P�dZ����P�M��@w���M�Q�M�5���E��   ��   �M���S���UR�M��5���}��uF�M��TF���E�P�M�Q�U�R��]�����M��_����uh���M��7h���E�P�M�J5���E�}�M�^2����tA�M���t$hd��M���Y���U���thl��M���g����E���th`��M��Y���M�Q�U�R�EP�q2�����E���MQj�UR��^�����E��]Ë�������������'���6���   










	�I ��Z�������������x������� 	
��T�4�t��� �I ����     ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�v^�����E]�����������U����D�����0  �D����A�E��D����D��}���   j�M���_���j$������   �U�����U��}���   �E����$�� j�\O����P�M��0V���   j�DO����P�M��V���|j�/O����P�M��V���gj�O����P�M���U���Rj�O����P�M���U���=j��N����P�M���U���(j��N����P�M��U���j��N����P�M��U���U�R�M��0���E� �j�M��^���E��j�M��^���E��]Ð	 ! 6 K ` � � u �  ���������������������������������������������������������������������������������������������������U���0  �M��XN���E� �D�����5  �   k� �D����$u8�EP�M�Q�UR�E�P�{'�����M���,����u�M�Q�M�/���E�  �D����A|	�E�A   ��E�   �D��+UԉU��M���M���M��M���E�   �E��E��}�t�}�tw�}���   �#  ��!����tZ�R_����tQ�M��L,����u2j	��L����P������Qj �U�R�M��OF�����U��P�M��]���j	�L����P�M��S����   �!����tQ�M���+����u2j�L����P������Pj �M�Q�M���E�����T��P�M������j�]L����P�M��1S���f�%!����tT�M��+����u5j
�3L����P��(���Rj ��x���P�M��E�����]T��P�M�����j
��K����P�M���R����E�    �}� ��   �D����D��   k� �D����$u8�EP�M�Q�UR�E�P�%�����M���*����u�M�Q�M�-���E�  �D����A|	�E�A   ��E�   �D��+UЉU��}� �����D����t�D����D��}��|  �EP�M���j���M�Q�U�R�M���E��P�M�����M��K*����u,�E�P��h���Qj �����R�M��RD������E��P�M��`���M��*����u,�E�P��X���Qj ������R�M��D�����E��P�M��(���E����  �} tj�M�Z���E�  �M���tw�E�PhT���H���Q�0����P�M������D����t,�M�Q�����R��8���P�A�������	E��P�M������M�Qj�U�R�.V����P�M�����!�D����t�U�R��@����P�M��p5���D����uj�M��yk���3�D���E̋D����D��}�@tj�M��Y���E�  �U����tR�U����Uȃ}�t�?�} tj�M�Y���E�q  �E�P�M�Q��p���R�#�������%D��P�M�����#�E�����u��`���Q�y#����P�M��4���U���t!�E�Ph����P���Q�.����P�M��p���U���t!�E�Ph����@���Q�.����P�M��G���} ��   �M��'������   �M�*V����u�M��'����t:�M�_T����t�UR�M�������EPj ��0���Q�O����P�M���k���@�UR�� ���Pj �����Q�URj �� ���P��N�������A�����C��P�M��k���*�M�L'����u�MQj ������R�N����P�M��k���M��(���E���t�M���N���M�Q�M��)���E��   �j�M��W���E�   �   �} ux�M��&����ul�M�U����u�M�&����t�URj�EP�S�����E�u�9�MQ�URj ������P�MQj������R�aS�������@�����B���E�:�8�} u%�M�Y&����u�EPj�MQ�(S�����E��j�M�)W���E��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E��aj �M��rE��P�E�P�M��eE��P�MQ��8�����E��]�������������������������U��� �EP�M��&���D���U��}� t�}�?tq�}�Xt��   �E�Pj�MQ�P�����E��   �D����D��M��#����th���M��c���E�   ��E�PhX��MQ��)�����E�w�D����D��E��aj �M��D��P�E�P�M�Q�U�R��7����P�M��|���E�P�MQ��=�����E�$�U�R�M��%���E��E�P�MQ�=�����E��]����������������������������������������������������������������������������U���h��'����tH�T�%�����T�j �M�Q�9�����T���    �T��E�P�M�D%���E��  ��  �D����?��  �D����D��   k� �D����?uS�   �� �D����?u=�U�R�������D����t�D����D���E�P�M�$���E�9  �M�Q�wD�����M������E��M��[���E��M��!����u�U�R�M�u$���E��  �D������   �D����@��   �M�Q�
9�����M��X!������   �X���tn�X� �E�P�M�Q�M���<��P�M��j���D����@t>�M�Q�8����P�M��G���U�R�E�PhT��M�Q�M���I�����<��P�M�����)�U�R�E�PhT��M�Q�M��I�����Z<��P�M������}� t�M��#���}� t�M�����M�� ����u�M���"����t�U�R�M�M#���E��   �   �D����t�D����@ut�D����t�D����D��#*����t:�}� u4�M�������u(�M��4A��P�M�Q�;0�����U�R�M��"���E�U��E�P�MQ�0�����E�>�j�M��P���E�-�+�D����tj�M�P���E��j�M�P���E��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   V�E�    �D����Qu�E����D����D��D����uj�M�lO���E�W  �R  �D����0��   �D����9��   �}� tG�D�� ��/��EЉUԋD����D��U�R�E�P�M��R��P�M�Q�U�R�q$�����E��4�D�� ��/��EȉŰD����D��U�R�E�P�M��_R���E��M��M�U�R�M� ���E�  �  �E�    �E�    �D����@��   �D����uj�M�eN���E�P  �W�D����A|7�D����P*�E؋Uܱ��`���ȋ�D����A���M؉u��j�M�N���E��   �D����D��e����D���U�D����D��}�@tj�M��M���E�   �M��tX�}� t&�U�R�E�P�M��@Q��P�M�Q�U�R�#�����E���E�P�M�Q�M��Q���E�U�U�E�P�M�P���E�V�T�}� t&�M�Q�U�R�M���P��P�E�P�M�Q�"�����E���U�R�E�P�M���P���E��M��M��U�R�M�����E^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�D����tw�D����_ui�D��Q��t[�D��H��_uM�D����D��D����D��D����A�U��D����D��}�vj�M��K���E��M��;���E��]�������������������������������������������U��j�EP��I�����E]�����������U���8�RP����t�f$����u	�E�   ��E�    �E��E�M��s;���D���U�D����D��M��M��}�Y��   �U�����$���D����D�hy��M�XZ���E�   h���M��kA���kh���M��\A���\h���M��MA���Mh���M��>A���>h���M��/A���/�yO���E�U�R�M)����Ph���E�P������P�M�����M��:���}� t�M�Q�M�����U�R�[����P�M��]���E�P�M����E��]ð���N ����������������������������������������������������������������������������������������������������������������������U��EP������E]�������������U����M��;9���D������   �D���E��M���0�M��}�wH�U��$��h,��M��\?���>h4��M��M?���/�-h<��M��<?���hD��M��-?���j�M�H���E�~�D���M�D����D��E�E��M���1�M��}�w/�U�����$���M�QhL��U�R�����P�M��v	���E�P�M����E��j�M�H���E��]Ë�����p�    ���������������������������������������������������������������������������������������������U���0�M��7���D����D��D���U��}�At�}�BtU�}�C��   �   �} u,�E����&u	�E� ���M����*u	�M����D����D��  �} tj�M��F���E�  �E� j>�M�����D����D��p  �U����D����D��U  �   k� �D����t�   �� �D����uj�M�dF���E�$  �} tj�M�LF���E�  �   k� �D����0���   �� �D���LЉM��D����D��}�v/j,�M������E�3�QP�M��I��P�U�R�M��0��P�M����j>�E�P�M���.��P�M�����D����$u�D����D��j^�M�Q�M��.��P�M������D����t�D����D��
j�M���V���M��%���U�R�M�0���E��M�n5���E��]���������������������������������������������������������������������������������������������������������������������������������������������������������������U���,j h`�j�U�����E��}� t�M��4���E���E�    �E��E�M�Q�U�R������EP�M�Qj �U�R�E�P�n�������[-������.��P�M��i���M�Q�M�����E��]���������������������������������������������������U����   �D����u�URj�EP�?�����E�/  �D����6|�D����9~ �D����_tj�M�tC���E��  �D����6�U��D����D��}�)u[�D����t2�D����=�M��D����D��}�|�}�~�E�������EPj�MQ��>�����E�y  ��}� |�}�~�E������}��uj�M��B���E�L  �M���2���UR�M�����E����  �M�QhT���X���R�
����P�M������D����t;�U�R��H���P�M�Q�)����Pj ��h���R��8��������,��P�M������E�Pj�M�Q�>����P�M��o���D����t1�D����@u�D����D��j�M��A���E�m  ��M�Qj�UR�=�����E�Q  �V����t��(���P��>����P�M�������M�Q�>����P�M������U���tY�����t8�E�P�M�Q�U�R�����Pj ��8���P��7��������+��P�M�������x���Q�^����P�M���������t&�U�R�E�P�M�Q��(�������+��P�M��Q����U�R�(����P�M��H���M������u(j)�E�P�M�Qj(�U�R�M7��������)��P�M����j h`�j�}�����E�}� t�M���0���E���E�    �E�E��M�Q�U�R�J1����j)�E�P��p���Q������Pj(��`���R��6�������v)��P�M��S����T����t�E���t�M�Q�M��S���;����t��P���R�����P�M��iS�����@���P������P�M��A���]����t��0���Q�?5����P�M��.S����� ���R�%5����P�M�����}� t�E�P�M��� ���j�M�?���E��M�Q�M�c���E��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�<�����E]�����������U��Q�M��M��0����t2���E���U���
�P�ҋ�]���������������������U����M��E��xu�   k������E���E� �E���]�����������������U��Q�M��E��@��]����������������U����M��E��x t�M��I�����E���E� �E���]��������������������U����M��E��H�U���J�P�҈E��E���u�M��Q�E���H�B�ЈE��E���]�����������������������������U����M��E��x t�M��Q�E��H�T��U���E� �E���]���������������U���j'�EPj �M�Q��:����Pj`�U�R�3�������%���E��]��������������������������U����M��E������E�} t�MQ�U���Ѓ���   ��   �} w�E   �M��Q;U��   �}   v3��   jh`�h  �������E�}� t�M��C���E���E�    �E��E��}� tA�M��y t�U��B�M���U��E��B��M��U��Q�E��M��H�   +U�E��P�3��!��M��Q+U�E��P�M��Q�E��H�D
��]� ������������������������������������������������������������������������U����D����u3���   ��   �D����0|8�D����9*�D����/�M��D����D��E��   �   �E�    �D����@tY�D����u3��o�7�D����A|$�D����P�U����D���T
��U������6�D����D�뚋D���U��D����D��}�@t�����E���]���������������������������������������������������������������������U���  �M���)���M���)���E�    �E�    �D���M��D����D��E��EЃ}�_��  �M���P.�$�4.�D����D�j�M�]9���E��  �M��)���M����   ��<���R�4����Pj<��l���P�/����P�M��L���M��b���ȃ�>u
j �M����j>�M�����} t�U��D����u�U�R�M�
���E�>  �D����D��D��M�j j ��,���R�P4����P�M�������E��D��M������u4�   k���D����1u�U�Rj~��\���P��.����P�M������M��N����u�M�Q�M��K���U�R�M�
���E�  �G  �   k���D��
��P�Q�M��.���   �E�   �   k���D����4�P�M��b.����  �D���U��D����D��M��Mԃ}�_��  �U����.�$��.�D����D�j�M�t7���E��  �   k���D������P�M���-���_  �   k���D������R�M�F���E�  �1  �   k���D��
����Q�M��cF���M�� ���U�R�M�����E�P  ��  jhd��E�P�M������M���-���M�Q�M����E�  �   k���D������P�M��E���E��  �   k���D������R�M���,��j j �����P������P�M������M��?����u�M��c%����tj�M�6���E�  �M�Q�UR�M�� ���E�s  �  �  �   k���D��
����Q�M��f,���   k� �D����uj�EP�M�����E�  �   k� �D����0�M�x�}�rj�M�{5���E��  �U���X�P�M���+���D���U��D����D��M��M�U��0�U�}��;  �E��$�D/j �M�Q��������U�R�EP�M�Q��L���Rj �����P�M��"�������������E�S  �  �M�Q�U�R�M��s��j,��|���P������Q�����������P�M��	H��j,��t���R��d���P�^���������P�M���G��j,��T���Q��D���R�6���������P�M��G��j)��4���Pj ��$���Q�v2�������^��P�M��G��j'�UR�M��G���E�  �;�E�P�MQ�M�����E�l  �!�D����D�j�M��3���E�I  ��  �   k���D��
����Q�M��A*����  �D���E��D����D��U��U؃}� t�}�0t!�N�D����D�j�M�`3���E��  j h���M�Q��������M��*���U�R�M����E�  j�M�3���E�  �,  �D���M��D����D��E��E�M��A�M�}�	��   �U���`/�$�X/�   k���D����(�R�M�B���E�  �   k���D��
��(�Q�M���A���D����?u7�����Q�b�����P�M���E���D����@u�D����D�������R��#����P�M��E��h���M���6���E�P�M�����E��j�M��1���E�n�j�M��1���E�]�j�M��1���E�L�}� t
�M��2���-�M��� ����u!�M�Qh��������R�����P�M�������E�P�M�t���E��]ÍI B&a&�'�'�'�'�- )(J(q(�(,)�(;)�)�)�+�,�- 	

�*�*�+�+�+�,-        ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E����E�P�MQ�UR�EP�o*�����E��]�����������������������U��Q�E��a�E�P�MQ�UR�EP�/*�����E��]�����������������������U���<�M�����D���M��}�B��  �U���,5�$�5�MQj�UR�)�����E�s  h`��M��#���M������u
j �M�����EP�M�������D����D��E����U�R�M��3���P�E�P�MQ������E�	  �   �� �D����$tC�   �� �D����u�URj�EP�_(�����E��  �j�M�],���E�  �D����D��D���E��}�T�i  �M����5�$�p5�D����D��MQ�UR�	�����E�U  �D����D�j�MQ�UR�6=�����E�.  �D����D��E��aj �M�����P�M�Q�UR�E�P�[����P�MQ� �����E��   ��   h`��M��"���M�z�����u
j �M��{���UR�M��?����D����D��E����M�Q�M�����P�U�R�EP������E�|�D����D�j�M�+���E�^�I�D����D�hl��M�S:���E�;�&�EPj�MQ�&�����E�"j�M�*���E��UR�EP�'������E��]ÍI �23�2�2�4 ��4�3�3�3S404�4�4�4 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����D�����  �} t]�D����XuO�D����D��M������th���M�8���E��   ��URhX��EP��������E��   �D����Yu%�D����D��MQ�UR��������E�   �EP�M�Q�������M�������t �U�Rh���E�P������P�M��N����*�M��%����t�M�Qh���U�R�[�����P�M��"����E�P�M�����E���MQj�UR�#�����E��]�����������������������������������������������������������������������������������U����D������   �D����6|�D����9~�D����_un�UR�M��y6���M������u$�M� �����u�M�>$����u�EP�M��E:���M�������u�MQ�M��-:���U�R�EP�`�����E�   �Nj �MQ�UR�EP�M�Q�J
�����U���*u	�E�   ��E�    �M�Q�U�R�EP�7�����E�m�kj�M��O&���MQ�M��+���M�D�����u�UR�M��9���M�,�����u"�M� �����u
j �M��!	���EP�M��g9���M�Q�M������E��]�����������������������������������������������������������������������������������������������������U��EP�MQ�UR�EP�"�����E]�����������������U����D�����  �D����_�  �D����D��D����A�E��D����D��}���   �M��"���{�������   hT��M��)��j�����P�M��)���}� tk�U��҃�#U��U�E�E��}�t�}�t�h���M��V)���h���M��G)���j�M�r$���E�U�M���#M��M�th���M��)���j)�M��_���U�R�M�#����E��j�M�*$���E���M�N���E��]�����������������������������������������������������������������������������������������������U��D����@u"�D����D��EP�M�#����E���MQ�UR�3������E]��������������������������U����   �M��x���E� �M���������  �D������  �D����@��  �X���t�Y���u�E�P�M������E�-  �M��������uH�M�QhT��U�R�B�����P�M��	����E���t"�M�Qj[��d���R�#����P�M�������E� �D����?�  �D����D��D���M��U���$�U��}�-��  �E���A�$�A�   �� �D����_um�   ��D����?uX�D����D��E�P�M�Qj j ��4���R����������P�M��+����D����@u�D����D��F�E�P�M�Qj'��T���R�E�P������Pj`�����Q��������
�����.��P�M��������  �D����D��E�P�M�Qj j��D���R������������P�M������  j@hD��M��"���E�Ph����t���Q������P�M��S����<�������u�U�R�<�������l  �D����D��M�Q��$���Rj]�E�Pj j�M�Q�f��������	�����R��P�M�������E��  �M�����D����D�j j�E�P������M��#����uE�M��b�����u+�M�Q�U�RhT��E�P�M��?������
��P�M��z�����M�Q�M��l����
j�M��	���M�������u�D����@�w����M������u<j]�M�Q�U�Rj[��|���P�R����������P�M������D����D��
j�M�����*�U�R��l���P��\���Q� �������+
��P�M�������.�U�R��L���Pj j��<���Q���������	��P�M������ ����D���E�}� t�}�@tW�W�M��)�����tj�M�����;�M�Q��,���RhT������Pj������������������	��P�M��#�����
j�M������M�Q�M�����E��]Ë�B>�>t=�>"?@ ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���@�M��K��j j�E�P�����P�M��M����M��	����uN�D����tA�D����@t4�U�R�E�PhT��M�Q�U�R�o������������Z��P�M�������D����@u�D����D��b�D����tj�M��~���J�M��p�����tj�M��f���2�U�R�E�PhT��M�Qj�M��<�����8��������P�M��s����U�R�M�����E��]�����������������������������������������������������������������������������U����D����uj�M����E�T�R�D����?u3�D����D�j �U�R�����Pj-�EP�������E��j �MQ������E��]����������������������������������������U��EP�N������E]�������������U��Q�M��M�� �����t�E��EP�MQ�U���M���	�B�Ћ�]� �������������������������U����M��M�������uX�} u*�M��e%�����Ej h`��EP�P������E��M��M�} t �U�E�L�Q�UR�M�����E�E��  ��} t�M� �E��]� ����������������������������������������������U��Q�M��E��xujh���MQ�UR��&������E��]� ��������������U��Q�M��E;Es�M�U��B��M���M�E��]� ��������������������U����M��E��x t�MQ�UR�E��H����E���M�M��E���]� �����������������������U����M��EP�MQ�U��B�M���I�B�ЉE��M�;Ms�UR�E�P�M��Q�E���H�B�����E���]� �������������������������U��Q�M��E��HQ�U��BP�MQ�UR�%������]� ���������������������U��� �EP�M���'���D���U��D����D��}�@u�D���U��D����D��}�_tj�M�,���E�   �D����D�j �U�R�H����j �E�P�:�����D����t�D����@t�D����D��աD����u�D����D�j�M����E��D����D��M�Q�M�s����E��]�������������������������������������������������������������������������������U��Q�E+E�E��M;M�~�U��U�EP�MQ�UR�'  ���EE��]������������������������U��   k� �D��
��?uR�   �� �D��
��$uj�MQ�c������E�;�$�D����D�j j �EP�4������E��j j�MQ������E]������������������������������������������������U���|���3ŉE��E��M��M���Y��M���������  �D������  �D����@��  �E� �M��t�E� ��E��D����0�E�x6�}�	0�D����D��U�R�E�P�@�����P�M���(���<  �D��MčM�����E� �D����$uT�D��Q��$uE�D��H��Wu�E��D����D��"�D��H��Vu�D����D�������D����Xu!�D����D�h���M��z���,  �D����$u?�   �� �D����$t)�D����D��E�P�������P�M��������   �D����?��   �E�P�L�����������tkj�M�Q�M�����U�R������P�\����EЃ}� t�E�P�M���
���.h���M�Q�U�Rh���E�P�����������P�M��Q����.h���M�Q�U�Rh���E�P�a�����������P�M��!�����M�����P�M�Q�{�����P�M������D�+Uă�~�@��J�����u�E�P�@��{����M�������u3�M��t
j,�M������U�R�M���&���E��thP�M�����0����Y� �M�Q�M�����E�M�3��������]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���  ���3ŉE��D���M��D����D��E���l�����l���T��  ��l������Q�$��Q�EP��������E��  �D����@u$�D����D�h���M�1!���E�  �3�����Q������P�URh����D����!�����:����E�t  �EP�v������E�`  ��T���Q�:�������\���R�+�������T������������   ��\�����������   jd�   �� �L�Q��T����9����uj�M����E��  �   �� �   k� �T��T��   k� �T���-u%�   ��   �� �T��T��   ���D�.��   �� �D�.��\���R�EPje������Q�U�R�����������������������E�W  �j�M�]���E�C  ��d���P������������tMj�M�Q��d����Q���U�R�����P�\�����p�����p��� t��p���P�M�f���E��  �M���Du5h���UR��d���Ph����,���Q�A�����������E�  �3h���UR��d���Ph�������Q������������E�m  �h  j j ��L���R����������P�/�������L���Q�M�1����E�/  j{��x��������U���t�����t���H|3��t���J~�(��<���P������P��x����f"��j,��x��������M��M��U���F�U��}�wu�E��$�4R��4���Q������P��x����"��j,��x���������$���R�o�����P��x�����!��j,��x������������P�G�����P��x�����!��j}�MQ��x��������E�<�:�M�w����E�-�+�D����D�j�M�$���E�j�M����E�M�3�������]Ë�yQ�M�MDNaO0NuP<PjQ�Q 																																																																						�I Q�P7QQ�P����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   �   k� �D��
��?u�   �� �D��
��$tj�M�����E�|  �D����D��8��U�<��E��@��M�M��}����h����r����<����g���U��8���h����<���<����@��M������M������E� �D����?u,�D����D��U�Rj�E�P�������P�M��x����jj�M�Q������P�M��]����M�������t�X��U���uj�E�P�������Pj<�M�Q�^����P�M��:���M������Ѓ�>u
j �M������j>�M�������E��t�D����t�D����D��M�8��U��<��E�@��M�Q�M�L����E��]������������������������������������������������������������������������������������������������������������������������U����E��aj�M�����P�E�P�M������P�MQ�p������E��]�������������������������U���(�D����tg�D����Zu'�D����D��M�����P�M�>����E�^�0j)�UR�E�P�������Ph���M�Q���������T����E�,�*j)�URj�E�Ph���M��r������������&����E��]������������������������������������������U���x�E�    �D����_u�U��� @  �U��D����D��D����A�  �D����Z�  �D����A�E�D����D��U��� �  �U��E��t�M���    �M���U��������U��}���  �E�% �  t�M���������   �M��U��U���E�%�����E��M��M��U���U�t�}�t@�}�tq�   �E�% �  t�M���?�����@�M���U���������   �U�E�E��r�M��� �  t�U���?����ʀ   �U���E�%����   �E��M��M��;�U��� �  t�E�%?����E���M��������M܋U܉U���E���  �E��k  �E���E؃}���   �M��$�`�U���������   �U��   �E�%����   �E��s�M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��MԋUԉUЋEЉE����E���  �E��  �  �D����$��  �E� �D����D��D���Ũ}�R�]  �E���H`�$� `�U����d���� �  �U��D  �E�%�g�� �  �E��/  �M����d���� �  �M��  �U����d���� �  �U��  �E�%���� |  �E���  �D��Q��Pu�D����D��D����D��D���Eȃ}�Q��   �M����`�$��`�D����D�����  �D����D��D����0|C�D����95�D���D��D
ѣD��^���E��M���   �M��E��-  ��E���  �7�D����D��(���	  �E���  �E���  �E���  �E���  ��  �E���  �D����D���  �E��D����D��D����0|�D����5~$�D����t	�E���  ��E���  �E��z  �D����0�EċM��� �  �M��U��� �  t�E�%����   �E��M��M���U��������U��E��E��M���t�U���������   �U���E�%����   �E��Mă�t�U���    �U���E�%�����E��Mă��M�t�}�t@�}�tr�   �U��� �  t�E�%?�����@�E���M���������   �M��U��U��s�E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��;�M��� �  t�U���?����U���E�%�����E��M��M���E���  �E��  ��E���  �E��  �D����D���  �D����0��  �D����8��  �D���U��D����D��M�������M��U��U��E���0�E��}��?  �M��$�a�U��� �  t�E�%����   �E��=�M��� �  t�U���������   �U��E��E���M��������M��U��U��E��E��M��M��U��� �  t�E�%?�����@�E���M���������   �M��U��U��  �E�% �  t�M���������   �M��;�U��� �  t�E�%����   �E��M��M���U��������U��E��E��M��M��U��U��E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��  �M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M��U��U��E��E��M��� �  t�U���?����U���E�%�����E��M��M��   �U��������� @  �U��l�E�%���� `  �E��Z�M���������    �M��F�U��������� h  �U��2�E�%���� p  �E�� �M��������� x  �M���E���  �E��H�C�D����9u�D����D��E���  ��D����t	�E���  ��E���  �E���]Ð<Y>Y�X>Y�X>Y�X[Z�[�Y�Y�Y�Y�Y2[�\ 																																																																					��Z]ZtZ�Z[ ��v]^�^7_]_K_q_�_�_����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�D���M��}� t)�}�At�0�D����D�h��M�,���E�j�M�����E�j�M�����E��]������������������������������������U��EP�MQ�(������E]���������U����EP�M��,���h��M��  ���M�Q�������P�M����j}�M��0����D����@u�D����D��U�R�M������E��]�����������������������������������U���@�EP�M������M��$������b  �D�����Q  �E�P�M�Qj �U�R�E�P������������������P�M�谻���M���������  �D����@��   h��M�������M���������   �D������   �D����@txj'�M�Q�U�R������Pj`�E�P�i�����������P�M��>���D����@u�D����D��M��)�����t�D����@th��M��[����Z����M��������t �D����u
j�M���
��j}�M��y����D����@u�D����D��'�M�������t�U�Rj�E�P������P�M��i����M�Q�M������E��]�������������������������������������������������������������������������������������������������������������������U���p���3ŉE��D����0�M�x5�}�	/�D����D��E�P�MQ�<��v����E�N  �I  �M��l����D����?utj �M�Q�������P�M��b����D���EȋD����D��}�@t7�D����D��D����t	�E�   ��E�   �U�R�M�������  jhX��D�P��  ����u�E�X��D����D��7jhp��D�R�  ����u�E�p��D����D���E�    �}� ��   �M�Q�������v�����twj�U�R�M��G����E�P�����P�\����E؃}� t�M�Q�M������:h���M��~���h���U�R�E�P�M�Q�U�R�I������������P�M��%
���:h���M��B���h���E�P�M�Q�U�R�E�P������������P�M���	���P�M��t0�D����@u"�M�����P�M�褷���D����D��j@hD��M�����P�M��{����U��t�<��ʹ����u�E�P�<�������M�Q�M������E�M�3�������]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��T�% @  ]������������������U��Q�M��E��@������]����������U��Q�M��E��@������]����������U����M��E��8 u	�E�   ��E�    �E���]�������������������������U����M��E��8	u	�E�   ��E�    �E���]�������������������������U��Q�M��E��@������]����������U��Q�M��E��@������]����������U��Q�M��E��@������]����������U����M��M��������u�E��H��	��t	�E�   ��E�    �E���]�����������������������U����M��M�������u�E��H��
��t	�E�   ��E�    �E���]�����������������������U��Q�M��E��@������]����������U����M��E��H������	�E�   ��E�    �E���]����������������U��Q�M��M��������t3���E���U���
��ҋ�]����������������������U��Q�M��E��@��]����������������U��Q�M��   ��]�����������������U����M��E��x t�M��I�+����E���E�    �E���]�����������������U��QV�M��E��x }.�M��Q�E���H��Ћ��M��Q�E���H�����M��q�U��B^��]�����������������������U��Q�M��E��@��]����������������U��j�hnd�    P���3�P�E�d�    ����uM�������E�    j �������j�������j�������j���x����E������} |�}}kE����   k����M�d�    Y��]�����������������������������������������������������U��Q�M��E��H��   �U��J��]��������������������U��Q�M��E��H�� @  �U��J��]��������������������U��Q�M��E��H��   �U��J��]��������������������U��Q�M��E��H��    �U��J��]��������������������U��Q�M��M�������u�E��H��   �U��J��]������������������������U��Q�M��E��H�� �  �U��J��]��������������������U��Q�M��E��H��   �U��J�E���]�����������������U��Q�M��E��@������]����������U��Q�E�    �	�E����E��M�;Ms�UU��EE���
�݋�]�����������������������������U��Q�E�    �	�E���E�M���t�E����E���E���]���������������U��} u3��G�E���Et.�M���t$�E��U�;�u�M���M�U���U�ǋE� �M�+�]���������������������������U��j�h�h�Ld�    P�ĜSVW���1E�3�P�E�d�    �} u3��   �E�    j���������u3��oj�ݴ�����E�    �EP�MQ�`������URj �EP�MQ�UR�M��p����M��:����E�`������E������   �j�������ËE�M�d�    Y_^[��]����������������������������������������������������������U��j�h0�h�Ld�    P�ĜSVW���1E�3�P�E�d�    �} u3��   �E�    j��������u3��pj�ͳ�����E�    �EP�MQ�`��|����U R�EP�MQ�UR�EP�M��_����M��)����E�`��
����E������   �j�������ËE�M�d�    Y_^[��]���������������������������������������������������������U��W�=@���   �}ww�U�����fn��p� ۹   #σ����+�3��of��ft�ft�f��#�uf��#���ǅ�EЃ������Sf��#���3�+�#�I#�[��ǅ�D�_���U��t93���   t�;�Dǅ�t G��   u�fn�f:cG�@�L�B�u�_�ø����#�f��ft �   #Ϻ������f��#�uf��ft@��f����t����뽋}3�������ك��E���8t3�����_�������������������������������������������������������������������������������������������U���0�E�E��M�Q�U��} t	�E�   ��E�    �E�E��}� u#h��hpjj j7h��j�?�������u̃}� u0�����    j j7h��h�h����������   �~  �} v	�E�   ��E�    �U�U�}� u#h�hpjj j8h��j�į������u̃}� u0�����    j j8h��h�h��g������   �  �   k� �E� �} ~�M�M���E�    �U��9Uv	�E�   ��E�    �E��E܃}� u#h �hpjj j=h��j� �������u̃}� u0�u���� "   j j=h��h�h ���������"   �_  �} t	�E�   ��E�    �U؉Uԃ}� u#h��hpjj j>h��j襮������u̃}� u0������    j j>h��h�h���H������   ��   �M��0�U����U��} ~A�E����t�U���EЋM����M���E�0   �U��EЈ�M����M��U���U빋E��  �} |>�M����5|3�E����E��M����9u�E�� 0�M����M���U�����M���U���1u�M�Q���E�P�&�M��Q���������P�U��R�EP�$�����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���@���3ŉE��E�    �E�    �EP�M��T����M�����Pj j j j �MQ�U�R�E�P������ �E�} t�M�UЉ�EP�M�Q�������E�U��u8�}�u�E�   �M��=����E��j��}�u�E�   �M��!����E��N�:�E��t�E�   �M������E��0��M��t�E�   �M�������E���E�    �M�������E܋M�3��t�����]��������������������������������������������������������������������U��j �EP�MQ�G�����]����������U���@���3ŉE��E�    �E�    �EP�M������M��4���Pj j j j �MQ�U�R�E�P�B����� �E�MQ�U�R�������E�E��u8�}�u�E�   �M�������E��j��}�u�E�   �M������E��N�:�M��t�E�   �M������E��0��U��t�E�   �M������E���E�    �M��o����E��M�3�������]������������������������������������������������������������������U��j �EP�MQ�d�����]����������U��j �EP�MQ�UR������]����������������������U��j �EP�MQ�:�����]����������U���@���3ŉE��E�    �E�    �EP�M��4����M�����Pj j j j�MQ�U�R�E�P������ �E�MQ�U�R�a������E�E��u8�}�u�E�   �M��+����E��j��}�u�E�   �M������E��N�:�M��t�E�   �M�������E��0��U��t�E�   �M�������E���E�    �M������E��M�3��b�����]������������������������������������������������������������������U��� �E�   �3�f�E��M�Q���  ��f�U��E�H�� �  f�M�U�B%�� �E�M��U��E��E�}� t�}��  t�P��  f�M��a�}� u)�}� u#�U�B    �E�     �Mf�U�f�Q�   �E�<  f�E��E�    ��M����  f�M��U����?  f�U��E���E�M�����U�B�E����M��U�B%   �uH�M���   �t	�E�   ��E�    �E�H��M��U�J�E���U�
f�E�f��f�E���M��U�ʋEf�H��]���������������������������������������������������������������������������������������������������U���,���3ŉE��EP�M�Q�������U�Rj j���ċM���U�Pf�M�f�H��������U�B�E֋M��UԋE�Pj jh��h �h8��M�Q�UR�EP������P�ް�����M�U�Q�E�M�3�������]������������������������������������������������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� ������������������������������������������������������SW3��D$�}G�T$���ڃ� �D$�T$�D$�}�T$���ڃ� �D$�T$�u�L$�D$3���D$���3�OyN�S�؋L$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$Oy���؃� _[� ���������������������������������������������̀�@s�� s����Ë�3������3�3������������������̀�@s�� s����Ë�3Ҁ����3�3�������������������U�� �]�������U���� ��E�M���u	�E�   ��E�    �U��U��}� u#h��hpjj j*h�j�4�������u̃}� u+�����    j j*h�hx�h����������E���M� ��E��]�������������������������������������������U����E%�����E�M#M��������   �} tj j �������U�3�t	�E�   ��E�    �M��M��}� u#h��hpjj j,h��j�L�������u̃}� u-�����    j j,h��hH�h����������   �/�} t�EP�MQ�������U���EP�MQ�k�����3���]��������������������������������������������������������������U��j�^�����]������������������S�܃������U�k�l$���   ���3ŉE��C���h�����h�����t����C���x�����x�������x�����x���wR��x����$��ǅ|���   �Cǅ|���   �7ǅ|���   �+ǅ|���   �ǅ|���   ��K�   ǅ|���    ��|��� ��   ��t����P�K��Q��|���R蕹������u{�C��p�����p���t��p���t��p���t� �M����M��U������U��C�@�]��	�M�����M��S��R�C��P�KQ��|���R��t���P�M�Q�e�����h��  ��t����P�������ǅl���    �K�9t�=P� u�SR腷������l�����l��� u�C�Q��������M�3�聾����]��[Ð����������ӄʄ����������������������������������������������������������������������������������������������������������������������������������������������U��3�]����������U��Q�E�    �E��U�+ȉM�u�M���t�E���E�M���M�σ}� }	�E�������}� ~�E�   �E���]����������������������������������U����E�E��M����tB�E�E��	�M����M��U����t�M���E��;�u
�E�+E����ыU����U�봋E�+E����]�����������������������������U��} u3��G�E���Et.�M���t$�E��U�;�u�M���M�U���U�ǋE� �M�+�]���������������������������U��Q�E���t=�U�U��	�E����E��M����t�E���U�;�u�E��֋M���M�3���]��������������������������������U���   ���3ŉE��E�H��  �U�JjU��P���P�k�������~Lj hj  h��h��h0���P���Q�a�������P��P���RjU�EP  P�Q�����P�h������M�3��L�����]��������������������������������������������U����E�Q���������u	�E�   ��E�    �U�E��B�M�QR���������u	�E�   ��E�    �E�M��H�U�z t	�E�   ��E�Q�D  ���E�U�E�Bj jh���3������M�Q��   t�E�H��   t�U�B��u
�M�A    ��]����������������������������������������������������������������U����E�Q���������u	�E�   ��E�    �U�E��B�M�y t	�E�   ��U�P�a   ���E��M�U��Qj jhP��P������E�H��u
�U�B    ��]�����������������������������������������U����E�    �} u3��X�Ef�f�M��U���U�E���A|	�M���Z~�U���a|'�E���z�M����M��Uf�f�E��M���M뾋E���]������������������������������U���   ���3ŉE��)����   ��x�����x����x tǅh���   �
ǅh���  j@��|���Q��h���R�EP蟗������u��x����A    �   ��  ��|���R��x����HQ貯�������  ��x����z tǅt���   �
ǅt���  j@��|���P��t���Q�UR�%�������u��x����@    �   �S  ��|���Q��x����P�9�������uf��x����Q��  ��x����Pj h�  h��h��h ��MQ�e�������P�URjU��x���P  P�U�����P�l������&  ��x����Q���  ��x����x ��   ��x����QR��|���P��x����R��������ua��x����H����x����Jj h�  h��h��h ��EP��������P�MQjU��x�����P  R詮����P��������}��x����H��uo�UR��  ����t_��x����H����x����Jj h�  h��h��h ��EP�;�������P�MQjU��x�����P  R�*�����P�A�������x����H��   ��   �f  ��x����z tǅl���   �
ǅl���  h�   ��|���P��l���Q�UR��������u��x����@    �   �4  ��|���Q��x����P����������  ��x����Q��   ��x����P��x����y ��   ��x����B   ��x����A�   k� ��x�����P  ��uJj h�  h��h��h ��EP��������P�MQjU��x�����P  R������P�������B  ��x����x ��   ��x����R賿������x���;A��   ��x���Rj�EP�a  ����t|��x����Q��   ��x����P�   k� ��x�����P  ��uJj h�  h��h��h ��UR�7�������P�EPjU��x�����P  Q�&�����P�=������{��x����B   ��x����A�   k� ��x�����P  ��uJj h�  h��h��h ��EP躾������P�MQjU��x�����P  R詫����P���������x����H��uǅp���   �
ǅp���    ��p����M�3��z�����]� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE��y����   �����������x tǅ���   �
ǅ���  jx�����Q�����R�EP��������u������A    �   �   �����R������Q��������u_j hL  h��h��h ��UR�G�������P�EPjU�������P  Q�6�����P�M�����������B��������A������B��uǅ ���   �
ǅ ���    �� ����M�3�������]� �������������������������������������������������������������������������������U��Q�} t�E���th���UR��������u5j�E�Ph  �M��P  Q芏������u3��^�}� u��P�Kh���UR�л������u'j�E�Ph   �M��P  Q�@�������u3����UR�������E��E���]�������������������������������������������������U������3ŉE�j	�E�PjY�MQ�̎������u3��j	�UR�E�P�&�������u�   �3��M�3��h�����]������������������������U��V�EP��������u,�} t&�M�R����������E�Q�������;�u3���   ^]�������������������������U����E�   �E�    �E�;Ed�}� t^�E�E�+����E�kM��U�
P�M�R�������E��}� ukE��M�T�E���}� }�M����M�	�U����U�딃}� u	�E�   ��E�    �E���]����������������������������������������������������U��������   �E��   k� 3ҋE�f��P  �M��A    �U�E���M���   �U��J�E��H���t�E���P�����Qh0��������U�����tw�U��B���t�U�R�j�������E�P�l������M��y uE�U�R�����Phh��i�������t'�M��Q���t�M�Q��������U�R��������E�P�@������M��y u3��  �} t�U��   �U���E�    �E�P�M�Q�E������E��}� t!�}���  t�}���  t�U�R� ��u3��G  �} t�E�M���} �*  �   k� 3ɋUf��   j h�   h��h �h8��E�P  P�>�������P�M���P  QjU�U��   R�*�����P�A�����j@�EPh  �M��   Q�E�������u3��   j@�U�   Rh  �E   P��������u3��vj_�M���   Q蓷������uj.�U�   R�{�������t'j@�E�   Pj�M��   Q���������u3��j
j�U��   R�E�P�w������   ��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���  ���3ŉE��	����   ��������������  ������MQ�  ��������������z tǅ ���   �
ǅ ���  h�   �����P�� ���Q�����R����u������     �   �   �����Q�������BP�l�������uD�����Q�  ����t1�����������B�����������Q��������������
��������uǅ����   �
ǅ����    �������M�3��w�����]� ������������������������������������������������������������������������������������U���膼���   �E��E��HQ�߳������u	�E�   ��E�    �U��E��Bjh�����M���u	�E�     ��]�����������������������������U��Q�E���  �U�
���E��E�M��H�U�E��B��]��������������U����ƻ���   �E��E��Q� �������u	�E�   ��E�    �U��E��B�M��QR��������u	�E�   ��E�    �E��M�H�U�B    �E��x t	�E�   ��M��R�M  ���E��E��M��Hjh�����U�%   t�M���   t
�E���u	�U�    ��]������������������������������������������������������������������U���覺���   �E��E��Q� �������u	�E�   ��E�    �U��E��B�M��y t	�E�   ��U��P�d   ���E�M��U�Qjh@����E���u	�U�    ��]��������������������������������������������������U����E�    �Ef�f�M��U���U�E���A|	�M���Z~�U���a|'�E���z�M����M��Uf�f�E��M���M뾋E���]����������������������������������������U���  ���3ŉE��I����   ������9������  ������MQ��  ���� ���������z tǅ����   �
ǅ����  h�   �����P������Q�� ���R����u������     �   ��  �����Q������BP謜��������  ������y tǅ����   �
ǅ����  h�   �����R������P�� ���Q����u������    �   �k  �����P������R�0�������u9��������  ������
������� ����H������� ����B��   ����������   ������x tu������QR�����P������R�ٷ������uO��������������
������� ����H������P�����������;Au������� ����B�B��������u5�� ���P�q  ����t"��������������������� ����Q��������   ��   ��  ������z tǅ����   �
ǅ����  h�   �����P������Q�� ���R����u������     �   ��  �����Q������P葚�������  ��������   ������������y t5������   ������������z u������� ����H�   ������z tj������Q�����������;BuN�����Pj�� ���Q�~  ����t0������   ������������z u������� ����H�0������   ������������z u������� ����H�   ������z uu������x ti�����Q������P�W�������uM�����Qj �� ���R��  ����t1��������   ������
������x u������� ����Q��������uǅ����   �
ǅ����    �������M�3��Y�����]� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���  ���3ŉE�艳���   �� ����y������  ������MQ�  ��������� ����z tǅ����   �
ǅ����  h�   �����P������Q�����R����u������     �   �$  �����Q�� ����P��������u^�� ����y u�����Rj�����P�Q  ����t1�����������Q�����������H���������������   �� ����z uu�� ����x ti�����Q�� ����P�[�������uM�����Qj �����R��  ����t1�����������H�����������B����������������������uǅ����   �
ǅ����    �������M�3��]�����]� ��������������������������������������������������������������������������������������������������������������������������U����E�    �Ef�f�M��U��U�E���E�}� tO�M���a|�U���f�E���'f�E���M���A|�U���F�E���f�E��M����U��DЉE�둋E���]����������������������������������������������U��Q�} t�E���th���UR誨������u0j�E�Ph  �M�QR����u3��Y�}� u��K�Fh���EP�e�������u"j�M�Qh   �U�BP����u3����MQ�y�����E��E���]�������������������������������������������U���f�Ef�E��E�    �	�M����M��}�
s�U��E��E��;�u3���ظ   ��]�������������������������U���V�E%�  �ȁ�   �щU��M����   �E�j�E�Ph   �M�Q����u3��9�U;U�t,�} t&�E��Q���������U��P�l�����;�u3���   ^��]������������������������������������������U����E�   �E�    �E�;Ed�}� t^�E�E�+����E�kM��U�
P�M�R�~������E��}� ukE��M�T�E���}� }�M����M�	�U����U�딃}� u	�E�   ��E�    �E���]����������������������������������������������������U���$���3ŉE��ܭ���   �E�jj �E�P薢����迭���  �E܋M܍U���E܋�M�} u�U�R�������(  �E�M��U�   �E�P�M�y t*�U�B���t�U��R�����Ph0��������M��    �U�: ��   �E������   �E�x t�M�Q���t�M�Q�1�������U�R�C������E�8 uO�M�Q�����Rhh���������t0�E�x t�M�Q���t�M�Q���������U�R��������0�E�x t�M�Q���t�M�Q���������U�R�Z������E�8 u3��!  �} t�M��   �M���E�    �U�R�E�P�������E�}� t!�}���  t�}���  t�M�Q� ��u3���   j�U�BP����u3��   �} t�M�U�jU�E�P  P�M�QR�������} txjU�E   P�M�QR������j@�EPh  �M�QR����u3��Cj@�E�   Ph  �M�QR����u3��j
j�E   P�M�Q�Բ�����   �M�3�躗����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E������E�    �E�    �} t	�E�   ��E�    �E؉Eԃ}� u#h��hpjj jmh�j�w������u̃}� u.������    j jmh�ht�h���K����������   �U�U��E����E��M��Q��U��E�    �E�    j �E�Pj@�MQ�UR�E�P�M�Q�b������E��E������   �Q�}� tJ�}� t8�U����E������P��T����E����M������P��T�M�Q�~t����Ã}� t�!����U܉�����E�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������U����E�    �E������E�E��M����M��U��B��E��E�    j �M�Q�U�R�EP�MQ�UR�|������E�}� t	�E�������E�E��E���]���������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�   ��E�    �E��E܃}� u&h��hpjj h�   h�j�#u������u̃}� u3�x����    j h�   h�h��h���ó�����   ��  �U������} t	�E�   ��E�    �E؉Eԃ}� u&h��hpjj h�   h�j�t������u̃}� u3�����    j h�   h�h��h���9������   �9  �} ��   �U�����u	�E�   ��E�    �EЉẼ}� u&h��hpjj h�   h�j�	t������u̃}� u3�^����    j h�   h�h��h��該�����   �   �E�    �UR�EP�MQ�UR�EP�MQ�U�R�ل�����E��E������   �[�}� tT�}� t@�E����U�������P��T����E����E� ������P��T�U�P��p����Ã}� t	�M������E�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    �E�P�MQ�u������u����8�U R�EP�MQ�UR�E�P�MQ�UR�v�����E�j�E�P讀�����E���]�������������������������������U��j�EP�MQ�UR�EP�MQ�\�����]��������������U��j �EP�MQ�UR�O�����]����������������������U���T�} u3���  �EP�M��/{���M������H�y u'�UR�EP�MQ莮�����EԍM��N����E��  �} t	�E�   ��E�    �U�U��}� u#h8�hpjj j>hX�j��p������u̃}� u=�B����    j j>hX�h��h8�萯�����E�����M��Ɗ���E��2  �} t	�E�   ��E�    �M�M�}� u#h��hpjj j?hX�j�ep������u̃}� u=躶���    j j?hX�h��h���������E�����M��>����E��  �E�EȋM���M�}� �  �Uf�f�E��M���M�M��
����P�E��L��t|�} u@3�f�U��M������@�M��D��t	�E�    �	�M��U�f�E�f�E��   �M���u	�E�    ��E����M�E��E���Ef�M�f�M��Uf�f�E��M���M�M��a����P�E��L��tM�} u3�f�U��?�E���E�M���u	�E�    ��E����M�E܋E���Ef�M�f�M��U��E�;�t/�M��U�;�~	�E�   ��E������E؉EčM��Ĉ���E��3�M���u�E�    �M�計���E���h����E�    �M�菈���E���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR襄����]����������������������U���XV�EP�M��+w���} u�E�    �M��e����E��	  �M��^����H�y u'�UR�EP�MQ蘧�����EЍM��-����E���  �} t	�E�   ��E�    �U�U��}� u#h8�hpjj j?h �j��l������u̃}� u=�!����    j j?h �hl�h8��o������E�����M�襆���E��I  �} t	�E�   ��E�    �M�M�}� u#h��hpjj j@h �j�Dl������u̃}� u=虲���    j j@h �hl�h���������E�����M������E���  �E�EċM���M�}� ��  �Uf�f�E��M���M�M������P�E��L���>  �} u@3�f�U��M�������@�M��D��t	�E�    �	�M��U�f�E�f�E���  �M���u3�f�E���   �M����U��f�M��M���M�u��M��Q����P�   k� �T
;�|C�u��M��1����@�   �� �T;�#�M������@�   ���T�E��f�E��b�u��M������H�   k��L;�|B�u��M��η���P�   ���L;�"�M�買���P�   k��T
�E��f�E��D�M�获���H�U��D��t�M��u����H�U���  �E���M��M�f�U�f�U��Ef�f�M��U���U�M��6����@�M��T���  �} u3�f�E��E  �M���M�U���u3�f�M���   �U����E��f�U��U���U�u��M��ʶ���@�   k� �D;�|C�u��M�誶���H�   �� �D;�#�M�莶���H�   ���D�M��f�M��b�u��M��g����P�   k��T
;�|B�u��M��G����@�   ���T;�"�M��+����@�   k��D�M��f�M��D�M������P�E��L��t�M������P�E���  �M���U��U�f�E�f�E��M��U�;�t/�E��M�;�~	�E�   ��E������U؉U��M�茂���E��3�E���u�E�    �M��p����E���Q����E�    �M��W����E�^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����Nk����teh��h@���P���E��}� u����c�E�   �E�E�M �M��E�    �U�U��E�    �E�P�MQ�UR�EP�MQ�U��#j �UU R�EP�MQ�UR�EP�MQ�T��]������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E������E�    �E�    �} t	�E�   ��E�    �E؉Eԃ}� u#h��hpjj jmh�j�e������u̃}� u.�ݫ���    j jmh�h��h���+����������   �U�U��E����E��M��Q��U��E�    �E�    j �E�Pj@�MQ�UR�E�P�M�Q�i�����E��E������   �Q�}� tJ�}� t8�U����E������P��T����E����M������P��T�M�Q�^b����Ã}� t�����U܉�����E�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������U����E�    �E������E�E��M����M��U��B��E��E�    j �M�Q�U�R�EP�MQ�UR蒘�����E�}� t	�E�������E�E��E���]���������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�   ��E�    �E��E܃}� u&h��hpjj h�   h�j�c������u̃}� u3�X����    j h�   h�h��h��裡�����   ��  �U������} t	�E�   ��E�    �E؉Eԃ}� u&h��hpjj h�   h�j�yb������u̃}� u3�Ψ���    j h�   h�h��h���������   �9  �} ��   �U�����u	�E�   ��E�    �EЉẼ}� u&h��hpjj h�   h�j��a������u̃}� u3�>����    j h�   h�h��h��艠�����   �   �E�    �UR�EP�MQ�UR�EP�MQ�U�R�%f�����E��E������   �[�}� tT�}� t@�E����U�������P��T����E����E� ������P��T�U�P��^����Ã}� t	�M������E�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   �E�    �E�    �E�    �E� �E�    ǅ`���   ǅd���    �E%�   tǅh���    �E��ǅh���   �E� j h:  h�h��h���M�Q������P�j�����U�� �  u/�E% @ t�M��ɀ   �M���}� �  t�U��ʀ   �U��E���E�t�}�t�}�t6�@�E�   ���   �M��t�U��   t	�E�   ���E�   @�   �E�   ��   �hd���     �E� ����3�t	�E�   ��E�    �U��U��}� u&h$�hpjj ha  h�j��^������u̃}� u3�!����    j ha  h�h��h$��l������   �  �M�M��U����U��}�pw_�E���D��$�,��E�    ��   �E�   ��   �E�   ��   �E�   �   �}�   �u	�E�   ��E�    �   �ac���     �U�����3�t	�E�   ��E�    �M���x�����x��� u&hh�hpjj h�  h�j�]������u̃�x��� u3�����    j h�  h�h��hh��\������   �   �E%   �E�}�   7�}�   tK�}�   �}�   t]�}� t3�}�   t6�d�}�   tO�Y�}�   t,�}�   t/�}�   t�<�E�   ��   �E�   ��   �E�   �   �E�   �   �E�   �   �!b���     �M�����3�tǅ|���   �
ǅ|���    ��|�����l�����l��� u&h$�hpjj h�  h�j�v\������u̃�l��� u3�Ȣ���    j h�  h�h��h$��������   �  �EȀ   �E�    �U��   t� ���#E%�   u�E�   �M��@t �U���   �U��E�   �E��M����M��U��   t�E�   �EȋM��    t�U���   �U��E�� t�M���   �M���U��t�E�   �E��Mw���M��U�:�u+�`���     �E� ����������    赡��� ��
  �M�   �U�R�E�P�M�Q��`���R�E�P�M�Q�UR�8������E�}���  �E�%   �=   ���   �M����   �U�������U��E�P�M�Q�U�R��`���P�M�Q�U�R�EP��������E�}��u^�M����E�������P��D
����M����M�	������P��D
��P�+Y����� ��� �E���	  �^�M����E�������P��D
����M����M�	������P��D
��P��X�����b���� �E��r	  �M�Q���E��}� ��   �E�    �U����M�������P��L����U����U�������P��L���E��M�Q�IX�����U�R���}� u�П���    �ş��� �E���  �}�u�M���@�M���}�u
�U����U��E�P�M�R�x�����E����E��M����E�������P��E��D
�M����E�������P��D
$$��M����M�	������P��D
$�E���H�  �M���   �  �U����   jj�j��E�Q������EЉUԋU�#Uԃ��u/�]���8�   t�E�Q�#�����谞����U���  �   3�f�E�j�M�Q�U�P�.x������uA�M���u8�U�R�E�P�M�R薍�������u�E�Q迈�����L�����U��\  j j j �E�Q� �����EЉUԋU�#Uԃ��u�E�Q�}������
�����U��  �E�%�   �  �M�� @ u'�U��� @ u�E @  �E��M��� @ M�M�U�� @ u&h��hpjj h�  h�j�.W������u̋M�� @ �M؁}�   &�}�   tW�}� @  t1�}�   t.�}� @ t%�D�}� @ t1�}�   t.�}� @ t%�'�E� �!�U��  ��  u�E��
�E���E��E%   �&  �E�    �E�    �E�    �M���@��  �U���   ��U��}�   @t'�}�   �t�}�   ���   �q  �E�   �e  �E�E��M����M��}���   �U��$���jj j �E�Q�>}������X�����\�����X����\���tPj j j �E�Q�}������@�����D�����@���#�D������u�E�Q聆����������U��  ��E�   �   �E�E��M����M��}���   �U��$���jj j �E�Q�|������H�����L�����H����L���tWj j j �E�Q�c|������P�����T�����P���#�T������u�E�Q�ԅ�����a�����U��q  �E�   ��E�   ��E�   �}� ��  j�E�P�M�R��t������p�����p��� ~7�}�u13�u&hL�hpjj h�  h�j�T������u��E�    ��p����U��}��t�}�t:�}�t"��   �E�Q������觚����U��  �}�﻿ u	�E���   �E�%��  =��  uO�M�R�܄����3�u&h��hpjj h  h�j��S������u��?����    �E�   �G  �U܁���  ����  uHj j j�E�Q��z�����EЉUԋU�#Uԃ��u�E�Q�W�����������U���  �E��Bj j j �E�Q�z�����EЉUԋU�#Uԃ��u�E�Q������蜙����U��  �}� ��   �E�    �E�    �E�    �E���t�����t���t��t���t��E���  �E�   ��E�﻿ �E�   �M�;M�~U�E�    �U�+U�R�EčL�Q�U�P�5x�����E��}��u�M�R�c���������� �E��   �M�M��M�룋U����M�������P��M����T$��
ыE����E� ������P��T$�U��   u	�E�    ��E�   �E����U�������P��U������D$$
M����M�	������P��D
$�E���HuH�M��t@�U����M�������P��L�� �U����U�������P��L�M���   ���   ���   �U����   �E�P���M�������M��E�   �U�R�E�P�M�Q��`���R�E�P�M�Q�UR�4������E�}��uk��P��O�����E����U�������P��T����E����E� ������P��T�U�P�
m����������M��"� �U����M�������P��M��E��]Ë�<�H�T�`�l��� �I �����������6�6���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�EP�MQ�UR�EP�MQ�R�����]��������������U���$�=4� ��  �E�    �} ��  �} t	�E�   ��E�    �E�E��}� u#h�hpjj jmh@�j�K������u̃}� u0�e����    j jmh@�h��h�賉���������D  �} t	�E�   ��E�    �U�U�}� u#h��hpjj jnh@�j�J������u̃}� u0�����    j jnh@�h��h���8�����������   �M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���M�U���U�E���Et�M���t�U��E�;��a����M��U�+ʉM܋E���j �EP�MQ�UR�z������]��������������������������������������������������������������������������������������������������������������������������U���4�E�    �} �@  �} t	�E�   ��E�    �E�E��}� u#h�hpjj j=h@�j�H������u̃}� u0�����    j j=h@�h��h��`�����������  �} t	�E�   ��E�    �U�U�}� u#h��hpjj j>h@�j�BH������u̃}� u0藎���    j j>h@�h��h�������������M  �MQ�M���Q���M�������   �����    ��   �M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���M�U���U�E���Et�M���t�U��E�;��a����i�M��U���P�M�R�kD����f�E��M��9���P�E�Q�OD����f�E��U���U�E���E�M���Mt�U���t�E��M�;�t��U��E�+ЉU܍M���`���E܋�]�������������������������������������������������������������������������������������������������������������������������������������������������������������������U���x  ���3ŉE�ǅ(���    ǅ����    ǅx���    ǅ����    ǅT���    ǅ���    ǅ4���    ǅ����    ǅ@���    �EP��`����bO��ǅ����    ǅp���    ǅ����    ǅ����    ǅ��������ǅ��������ǅ|�������ǅ��������ǅ��������ǅH���    蔋���������} tǅ����   �
ǅ����    ������������������ u&h�hpjj h  hx�j��D������u̃����� uI�)����    j h  hx�h��h��t�����ǅx���������`����^����x����1;  �E�������������Q��@��   ������P�w������\�����\����t-��\����t$��\�������\��������P��������
ǅ������������H$�����х�uV��\����t-��\����t$��\�������\��������P��������
ǅ������������B$�� ���ȅ�tǅ����    �
ǅ����   ������������������ u&hh�hpjj h	  hx�j�ZC������u̃����� uI謉���    j h	  hx�h��hh��������ǅ����������`����']���������9  �} tǅ����   �
ǅ����    ������������������ u&h��hpjj h  hx�j�B������u̃����� uI�����    j h  hx�h��h���N�����ǅ����������`����~\���������9  ǅ����    �E������ǅ����    �����������������������8  ������u������ u�8  ǅ����    ǅX���    ǅH���    ǅ ���    ǅ��������ǅx���    ǅ����    �������Uǅ��������ǅ|�������ǅ��������ǅ���������E��������������������E���E������ �5  ������ ��4  �������� |%��������x��������(����������
ǅ����    ������������k�����	��X�����H�����X�����X�����  �E���%��  �������u\j
��p���R�EP�1k������~9��p������$u+������ uh@  j ������P�g����ǅ����   �
ǅ����    �������.  j
��p���Q�UR��j��������������p������E������ ��   ������ |#��p������$u������d}ǅ����   �
ǅ����    ������������������ u&h�hpjj hU  hx�j��?������u̃����� uI�����    j hU  hx�h��h��]~����ǅ����������`����Y���������6  ������;�����~��������������������������������������   ��X�����   3�tǅ����   �
ǅ����    ������������������ u&h��hpjj ha  hx�j��>������u̃����� uI�%����    j ha  hx�h��h���p}����ǅ����������`����X���������-5  ��X����������������2  �������$�d������ u	������t������u�������u��1  ǅ@���    ��`����:���P������R�I���������   ������P�MQ������R�#I  ���E��������U���U��������tǅ����   �
ǅ����    ������������������ u&h�hpjj h�  hx�j�y=������u̃����� uI�˃���    j h�  hx�h��h��|����ǅ����������`����FW����������3  ������P�MQ������R�FH  ���0  ǅ���    �������4�����4�����x�����x�����T���ǅ����    ǅ��������ǅ@���    �O0  ��������$�����$����� ��$�����$���wj��$�������$�����������������E���������������4���������������#�������ɀ   ����������������������/  ��������*��  ������ u�MQ��R������x����  j
��p���R�EP�Rf��������|�����p������M������ �'  ��|��� |#��p������$u������d}ǅ����   �
ǅ����    ������������������ u&h �hpjj h�  hx�j�J;������u̃����� uI蜁���    j h�  hx�h��h ���y����ǅp���������`����U����p����1  ��|���;�����~��|������������������������������������|����������� uE��|�����Ǆ����   ��|�������������������|�������������������   ������Q������Rj��|�����������Q�l������tǅ����   �
ǅ����    ������������������ u&h��hpjj h�  hx�j��9������u̃����� uI�?����    j h�  hx�h��h���x����ǅ����������`����S���������G0  �/-  �+��|�������������h�����h���P�MP������x�����x��� }����������������x����ډ�x����k�x���
�������TЉ�x����,  ǅ����    �,  ��������*��  ������ u�MQ��O�����������  j
��p���R�EP�Ec��������������p������M������ �'  ������ |#��p������$u������d}ǅ���   �
ǅ���    ����������������� u&h��hpjj h�  hx�j�=8������u̃����� uI�~���    j h�  hx�h��h����v����ǅ����������`����
R���������.  ������;�����~��������������������������������������������������� uE��������Ǆ����   ������������������������������������������   ������Q������Rj��������������Q�i������tǅ����   �
ǅ����    ���������������� u&h8�hpjj h�  hx�j��6������u̃���� uI�2}���    j h�  hx�h��h8��}u����ǅ`���������`����P����`����:-  �"*  �+��������������������������P�@M���������������� }
ǅ���������k�����
�������DЉ�������)  ������������������I����������.�B  ���������$���U���lu�M���M��������   �����������������������   �M���6u+�E�H��4u�U���U������ �  �������   �M���3u(�E�H��2u�U���U������%����������e�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu��������   �������ǅX���    �����"�������� �������������   �������S(  �������� ����� �����A�� ����� ���7��%  �� �����0�$����������0  u������   ��������������  ��  ǅt���    ������ u�UR�mp����f��,����  ������ |������d}ǅ����   �
ǅ����    ������������������ u&h��hpjj h�  hx�j�3������u̃����� uI�z���    j h�  hx�h��h���[r����ǅX���������`����M����X����*  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R�d������tǅ|���   �
ǅ|���    ��|��������������� u&h@�hpjj h�  hx�j�2������u̃����� uI��x���    j h�  hx�h��h@��%q����ǅ����������`����UL����������(  � #  �,����������������P�����P���Q�Jn����f��,�����,���Rh   ������P������Q�ty������t�����t��� t
ǅ4���   �^  ������ u�UR�H����f��8����  ������ |������d}ǅ����   �
ǅ����    ��������l�����l��� u&h��hpjj h�  hx�j�>1������u̃�l��� uI�w���    j h�  hx�h��h����o����ǅ����������`����K���������'  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R�4b������tǅ����   �
ǅ����    ��������d�����d��� u&h��hpjj h�  hx�j�0������u̃�d��� uI�Zv���    j h�  hx�h��h���n����ǅH���������`�����I����H����b&  �   �,��������������������������Q�hF����f��8����   k� ��8���������ǅ����   �������������B   ������ u�EP�F������D����  ������ |������d}ǅ����   �
ǅ����    ��������\�����\��� u&h��hpjj h�  hx�j��.������u̃�\��� uI�"u���    j h�  hx�h��h���mm����ǅ@���������`����H����@����*%  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������P������Qj��������������P��_������tǅ����   �
ǅ����    ��������T�����T��� u&h��hpjj h�  hx�j�-������u̃�T��� uI��s���    j h�  hx�h��h���7l����ǅ����������`����gG����������#  �2  �+����������������8�����8���R��C������D�����D��� t��D����x u#�p�������������R�W�����������d������%   t/��D����Q��������D���� �+���������ǅ@���   �(ǅ@���    ��D����Q��������D�����������d  ��������0  u������   �������������uǅ����������������������������<��������� u�EP��B�����������  ������ |������d}ǅL���   �
ǅL���    ��L��������������� u&h��hpjj h:  hx�j�+������u̃����� uI��q���    j h:  hx�h��h���Cj����ǅ����������`����sE��������� "  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������P������Qj��������������P�\������tǅD���   �
ǅD���    ��D��������������� u&h��hpjj h>  hx�j�p*������u̃����� uI��p���    j h>  hx�h��h���i����ǅ0���������`����=D����0�����   �  �+��������������������������R��@����������������%  ��   ������ u�t�������ǅ@���   �������������<�����(�����<�������<�����(��� t��������t������������뾋����+��������������t������ u�p��������������������<�����������<�������<��������� t��������t������������뾋����+�������������  ������ u�UR�?�����������  ������ |������d}ǅ<���   �
ǅ<���    ��<��������������� u&h��hpjj h�  hx�j�\(������u̃����� uI�n���    j h�  hx�h��h����f����ǅ ���������`����)B���� ����  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R�RY������tǅ4���   �
ǅ4���    ��4��������������� u&h��hpjj h�  hx�j�&'������u̃����� uI�xm���    j h�  hx�h��h����e����ǅ����������`�����@���������  �  �+������������������������Q�=�����������R^������   3�tǅ,���   �
ǅ,���    ��,��������������� u&h�hpjj h�  hx�j�@&������u̃����� uI�l���    j h�  hx�h��h���d����ǅ����������`����@���������  ��  �������� t������f������f���������������ǅ4���   �  ǅ���   �������� ��������������@��������������  ������ ��  ������ |������d}ǅ$���   �
ǅ$���    ��$��������������� u&h��hpjj h�  hx�j�	%������u̃����� uI�[k���    j h�  hx�h��h���c����ǅ���������`�����>��������c  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R�V������tǅ���   �
ǅ���    ����������������� u&h(�hpjj h�  hx�j��#������u̃����� uI�2j���    j h�  hx�h��h(��}b����ǅ����������`����=���������:  �x  ������������ǅ ���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Yh�  hp�j��������]  Q�������H�����H��� t��H���������������]  �� ����
ǅ�����   ������ u#�M���M�U�B��J���|����������!  ������ |������d}ǅ���   �
ǅ���    ����������������� u&h��hpjj h  hx�j�3"������u̃����� uI�h���    j h  hx�h��h����`����ǅ���������`���� <��������  ������t&h��hpjj h  hx�j�!������u̋������������������������������������B��J���|�����������`����n��P�����R������P������Q�� ���R������P��|���Q�   k���0�Q��Ѓ���������   t6������ u-��`����n��P������P�   k�	��0�P��Ѓ���������gu;��������   u-��`�����m��P������P�   ����0�R��Ѓ����������-u!��������   ��������������������������Q�{J�����������?  ��������@������ǅ0���
   �   ǅ0���
   �   ǅ����   ǅ(���   �
ǅ(���'   ǅ0���   ������%�   t2�   k� Ƅt���0��(�����Q�   �� ��t���ǅT���   �)ǅ0���   ��������   t������   �������������� �  �N  ������ u�UR�yN�����������������#  ������ |������d}ǅ����   �
ǅ����    ������������������ u&h��hpjj h�  hx�j��������u̃����� uI�Fe���    j h�  hx�h��h���]����ǅ����������`�����8���������N  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R��O������tǅ����   �
ǅ����    ������������������ u&h�hpjj h�  hx�j�������u̃����� uI�d���    j h�  hx�h��h��[\����ǅ ���������`����7���� ����  �V  �1����������������t�����t���Q�QL������������������  ��������   �N  ������ u�EP�L�����������������#  ������ |������d}ǅ����   �
ǅ����    ��������x�����x��� u&h��hpjj h�  hx�j�������u̃�x��� uI��b���    j h�  hx�h��h���1[����ǅl���������`����a6����l�����  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������P������Qj��������������P�M������tǅp���   �
ǅp���    ��p�����h�����h��� u&h��hpjj h�  hx�j�^������u̃�h��� uI�a���    j h�  hx�h��h����Y����ǅd���������`����+5����d����  ��  �1����������������\�����\���R��I�����������������r	  �������� ��  ��������@�R  ������ u�UR�z1�������������������%  ������ |������d}ǅ`���   �
ǅ`���    ��`�����X�����X��� u&h��hpjj h�  hx�j�&������u̃�X��� uI�x`���    j h�  hx�h��h����X����ǅT���������`�����3����T����  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R�K������tǅP���   �
ǅP���    ��P�����H�����H��� u&h��hpjj h�  hx�j��������u̃�H��� uI�B_���    j h�  hx�h��h���W����ǅL���������`����2����L����J  �	  �3����������������D�����D���Q�P/�������������������Q  ������ u!�UR�(/��������������������'  ������ |������d}ǅ@���   �
ǅ@���    ��@�����8�����8��� u&h��hpjj h�  hx�j��������u̃�8��� uI�$^���    j h�  hx�h��h���oV����ǅ<���������`����1����<����,  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R��H������tǅ0���   �
ǅ0���    ��0�����(�����(��� u&h��hpjj h  hx�j�������u̃�(��� uI��\���    j h  hx�h��h���9U����ǅ4���������`����i0����4�����  �4  �5����������������,�����,���Q��,��������������������  ��������@�P  ������ u�EP��,������������������$  ������ |������d}ǅ ���   �
ǅ ���    �� ������������� u&h��hpjj h  hx�j�p������u̃���� uI��[���    j h  hx�h��h���T����ǅ$���������`����=/����$�����  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������P������Qj��������������P�fF������tǅ���   �
ǅ���    ��������������� u&h��hpjj h  hx�j�:������u̃���� uI�Z���    j h  hx�h��h����R����ǅ���������`����.��������
  ��  �2������������������������R�*������������������M  ������ u�EP�s*����3ɉ������������%  ������ |������d}ǅ ���   �
ǅ ���    �� ��������������� u&h��hpjj h4  hx�j�������u̃����� uI�qY���    j h4  hx�h��h���Q����ǅ���������`�����,��������y	  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������Q������Rj��������������Q�D������tǅ����   �
ǅ����    ������������������ u&h��hpjj h8  hx�j��������u̃����� uI�;X���    j h8  hx�h��h���P����ǅ���������`����+��������C  �  �3��������������������������P�I(����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�L�����P�����������   ���������������L�����������P����������� �  u(������%   u��L�����P����� ��L�����P��������� }ǅ����   �%���������������������   ~
ǅ����   ��L����P���u
ǅT���    �   i��  �������������������������������������������� ��L����P�����   ��0����RP��P���R��L���P�)����0�������0����RP��P���Q��L���R��'����L�����P��������9~������(�����������������������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0��������������������u������ u�  ��4��� �b  ��������@tv��������   t�   k� Ƅt���-ǅT���   �L��������t�   k� Ƅt���+ǅT���   �%��������t�   k� Ƅt��� ǅT���   ��x���+�����+�T�����������������u������Q�UR������Pj �7  ��������Q������R�EP��T���Q��t���R�_  ����������t'��������u������R�EP������Qj0��  ����@��� ��   ������ ��   ǅ����    �������������������������������������������������������� ��   ������f�f������������Rj�E�P������Q��T������������������������������ u	������ uǅ���������*������P������Q�UR������P�M�Q�D  ���N����(������R������P�MQ������R������P�  �������� |'��������t������R�EP������Qj �  ����H��� tj��H���R�����ǅH���    �������X��� t��X���tǅ����    �
ǅ����   ������������������ u&hh�hpjj h�  hx�j��������u̃����� uI�QR���    j h�  hx�h��hh��J����ǅ����������`�����%���������Y  �������*  ������ �  ǅ����    ���������������������;�������  �������������������������������������  ������$�h���������E�������MQ��!�����  ���������E�������MQ�$G�����d  ���������E�������MQ�!�����@  ���������E�������MQ�9�����  ���������E�������MQ�9������   ���������E�������MQ�2!������   ���������E�������MQ�DY�����������������   3�tǅ����   �
ǅ����    ������������������ u&h��hpjj h2	  hx�j��	������u̃����� uF�P���    j h2	  hx�h��h���gH����ǅ����������`����#���������'������1�����������������`����n#���������M�3��(����]ÐN��������������N�_�=�,�s��� �I ���������� ���,�4��V� K�Y����S�w��   	
����6�Z����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���<�E�    �E�    �E�H��pt	�U��pu'�E�H�U;�u	�E�   ��E�    �E��  �E�H��st�U�B��St	�E�    ��E�   �M��M��U��st�E��St	�E�    ��E�   �M�M��}� u�}� ta�U�;U�uJ�E�H��  t	�E�   ��E�    �U��  t	�E�   ��E�    �E�;E�u	�E�   ��E�    �E���  �M�Q��dtv�E�H��itj�U�B��ot^�M�Q��utR�E�H��xtF�U�B��Xt:�M��dt1�U��it(�E��ot�M��ut�U��xt�E��X�,  �M�Q��dtE�E�H��it9�U�B��ot-�M�Q��ut!�E�H��xt�U�B��Xt	�E�    ��E�   �M��dt6�U��it-�E��ot$�M��ut�U��xt�E��Xt	�E�    ��E�   �M�;M�t3��   �U�B%   t	�E�   ��E�    �M��   t	�E�   ��E�    �U�;U�u;�E�H�� t	�E�   ��E�    �U�� t	�E�   ��E�    �E�;E�t3���M�;Uu	�E�   ��E�    �Eċ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E����U�
�E��A��Q�]��������������������U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�3�����E��}��u�M�������U����M���]�������������������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��|�U�    �E�E��M���M�}� ~N�U��E��MQ�UR�E�P�w������M���M�U�:�u�E�8*u�MQ�URj?�L�������띋E�8 u�M�U���]������������������������������������������������U���P  ���3ŉE�ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    �EP��P�������ǅ����    �8����p����} tǅD���   �
ǅD���    ��D������������� u&h�hpjj h  hx�j���������u̃���� uI�38���    j h  hx�h��h��~0����ǅ����������P�������������  �E�� ����� ����Q��@��   �� ���P��$�����������������t-�������t$�������������������P��������
ǅ������������H$�����х�uV�������t-�������t$�������������������P��������
ǅ������������B$�� ���ȅ�tǅL���    �
ǅL���   ��L������������� u&hh�hpjj h	  hx�j�d�������u̃���� uI�6���    j h	  hx�h��hh��/����ǅ����������P����1
���������A  �} tǅ���   �
ǅ���    �������<�����<��� u&h��hpjj h  hx�j��������u̃�<��� uI�6���    j h  hx�h��h���X.����ǅ����������P����	���������  ǅ����    ǅ����    ǅ����    ǅ����    ǅ|���    �E��������������������E���E������ �i  ������ �\  �������� |%��������x��������(���������
ǅ���    �����������k�����	��������H�����������������   3�tǅ4���   �
ǅ4���    ��4��������������� u&h��hpjj he  hx�j�5�������u̃����� uI�4���    j he  hx�h��h����,����ǅ����������P�������������  ��������,�����,����%  ��,����$��Iǅ����    ��P�����:��P������R��;��������   ������P�MQ������R�  ���E��������U���U��������tǅ���   �
ǅ���    �������$�����$��� u&h�hpjj h�  hx�j��������u̃�$��� uI�V3���    j h�  hx�h��h��+����ǅ����������P���������������  ������P�MQ������R��  ����  ǅ����    ������������������������������������ǅ����    ǅ��������ǅ����    �  �������������������� ������������wj�������� J�$�J���������������E���������������4���������������#�������ɀ   ����������������������  ��������*u:�MQ�s���������������� }���������������������؉������k�����
�������DЉ������  ǅ����    �  ��������*u'�UR����������������� }
ǅ���������k�����
�������TЉ������F  ��������������������I������������.�3  ��������HJ�$�4J�M���lu�E���E��������   �����������������������   �E���6u,�U�B��4u �M���M�������� �  �������   �E���3u)�U�B��2u�M���M������������������S�E���dt7�U���it,�M���ot!�E���ut�U���xt�M���Xu�ǅ����    ������#�������� ���������������   ��������  ��������������������A������������7�)
  ���������J�$�xJ������%0  u��������   ��������������  t[ǅ����    �EP�J%����f��t�����t���Qh   ������R������P�t0���������������� t
ǅ����   �2�MQ������f��l����   k� ��l���������ǅ����   �������������J	  �EP�T����������������� t�������y u#�p�������������P�`�����������e��������   t/�������B��������������+���������ǅ����   �(ǅ����    �������B��������������������  ������%0  u��������   �������������uǅ������������������������������MQ�T�������������������  ��   ������ u�t�������ǅ����   �������������������������������������������� t���������t��������������뾋�����+��������������u������ u�p��������������������������������������������������� t���������t��������������뾋�����+������������*  �MQ�4�������8���� ������   3�tǅH���   �
ǅH���    ��H�����@�����@��� u&h�hpjj h�  hx�j���������u̃�@��� uI�@,���    j h�  hx�h��h��$����ǅ����������P���������������	  �_  �������� t��8���f������f����8����������ǅ����   �%  ǅ����   �������� ��������������@������������������ǅ|���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Zh�  hp�j��������]  R������������������ t ��������������������]  ��|����
ǅ�����   �U���U�E�H��P���������������P����`1��P������P������Q������R��|���P������Q������R�   k���0�R��Ѓ�������%�   t6������ u-��P�����0��P������Q�   k�	��0�Q��Ѓ���������gu:������%�   u-��P����0��P������Q�   ����0�P��Ѓ����������-u ������   ��������������������������R�W������������  ��������@������ǅ����
   �   ǅ����
   �   ǅ����   ǅ����   �
ǅ����'   ǅ����   ��������   t2�   k� Ƅ����0��������Q�   �� ������ǅ����   �)ǅ����   ������%�   t��������   �������������� �  t�EP�a�����������������   ��������   t�UR�6�����������������   �������� tE��������@t�UR�����������������������EP����������������������@��������@t�UR���������������������EP�p�����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ������������������ }ǅ����   �%���������������������   ~
ǅ����   �����������u
ǅ����    �   i��  �������������������������������������������� �������������   �������RP������R������P������0�������������RP������Q������R�����������������������9~���������������������������������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0�������������������� �b  ��������@tv��������   t�   k� Ƅ����-ǅ����   �L��������t�   k� Ƅ����+ǅ����   �%��������t�   k� Ƅ���� ǅ����   ������+�����+�������`�����������u������Q�UR��`���Pj �
  ����p���Q������R�EP������Q������R�
  ����������t'��������u������R�EP��`���Qj0�+
  �������� ��   ������ ��   ǅ0���    ��������h�����������d�����d�����������d�������d��������� ��   ��h���f�f��z�����z���Rj�E�P��(���Q�%������0�����h�������h�����0��� u	��(��� uǅ���������*��p���P������Q�UR��(���P�M�Q�	  ���N����(��p���R������P�MQ������R������P�c	  �������� |'��������t������R�EP��`���Qj ��  �������� tj������R�O�����ǅ����    �i��������� t������tǅ ���    �
ǅ ���   �� ������������� u&hh�hpjj h�  hx�j�=�������u̃���� uF�"���    j h�  hx�h��hh�������ǅ����������P����
������������������������P���������������M�3�������]Ë��79h9�9_:n:�:<�9�9�9�9�9�9 �I 7;�;�:<< �L@\<�=�B'=f@{<}BG?C�B�=�B�BqF   	
����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP������E��}��u�M�������U����M���]�������������������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��|�U�    �E�E��M���M�}� ~N�U��E��MQ�UR�E�P�w������M���M�U�:�u�E�8*u�MQ�URj?�L�������띋E�8 u�M�U���]������������������������������������������������U��Q�����9(�u	�E�   ��E�    �E���]����������������������U��Q�E�E��M�Q�UR�EP���������]���������������U��Q�E�E��M�Qj �UR���������]�����������������U��Q�E�E��M�Q�UR�EP��������]���������������U��Q�E�E��M�Q�UR�EP�e�������]���������������U��������9(�u	�E�   ��E�    �M��M�} t������U���E�    �E��(��E��]���������������������������U��j�h �h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h��hpjj j6h��j���������u̃}� u.�"���    j j6h��h0�h���p��������   �U�U��k���    �� �Pj�������E�    �J���    �� �P��������EԋE�Pj �MQ�%���    �� �P�L�����E��
���    �� �P�U�R�O�����E������   ������    �� �Pj�����ËE܋M�d�    Y_^[��]������������������������������������������������������������������������������������������������U��Q�E�E��M�Qj �UR���������]�����������������U��� �E������EP�M�������M��E��P�MQ�M��7����BtP�MQ�U�R�������E�}� u�E��E���E������M��M��M�������E���]�������������������������������U���H�} u�} v�} t	�E�     3��  �} t	�M������}���w	�E�   ��E�    �U��U�}� u#h@�hpjj jJhx�j�:�������u̃}� u0����    j jJhx�h��h@��������   �  �MQ�M������M������   �����    �  �M���   ~C�} t�} v�URj �EP�������
��� *   ������M܍M������E��  �} ��   �} v	�E�   ��E�    �U��U�}� u#h�hpjj j]hx�j�;�������u̃}� u=���� "   j j]hx�h��h��������E�"   �M������E��}  �M�U��} t	�E�    �E�    �M�������E��O  �B  �E�    �M�Qj �UR�EPj�MQj �M������BP��E��}� t
�}� ��   �}� ��   ����z��   �} t�} v�MQj �UR�T�����3�t	�E�   ��E�    �M�M��}� u#h��hpjj j{hx�j��������u̃}� u:�\��� "   j j{hx�h��h���
�����E�"   �M�������E��L�"��� *   ���� �E̍M������E��*�} t�M�U���E�    �M������E���M�������]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�����j �EP���P�MQ�U�R�������E�}� u�E��E���E������E���]������������������������U��j �EP�MQ�UR�EP������]�����������������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� �������������������������������������������U���$�E=��  u	f�E�)  �MQ�M������M��X����   �����    u>�M��A|�U��Z�E�� �E���M�M�f�U�f�U��M�����f�E���   �E=   }Yj�MQ��������uf�Uf�U��M������f�E��   �+�M������ �M���   f�
f�E��M�����f�E��`j�M�Qj�URh   �M����� �   �ዔ�   R�n������uf�Ef�E��M��T���f�E��f�M�f�M�M��>���f�E��]������������������������������������������������������������������������������������������U��j �EP�������]�������������U��j
j �EP������]������������U��EPj
j �MQ�����]��������U��EP�MQ������]������������U��EPj
j �MQ�������]��������U��EPj
j �MQ�����]��������U��EP�����]����������������U��j
j �EP�K�����]������������U��j
j �EP������]������������U��j j j�EP�MQ�UR�O����]������������������U��j�h �h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j�,������E�    �EP�MQ�UR�EP�MQ�UR�[   ���E��E������   �j�C�����ËE�M�d�    Y_^[��]����������������������������������������U����} t	�E�   ��E�    �E�E��}� u&h� hpjj hX  h �j�k�������u̃}� u3�����    j hX  h �hh� ������   �G  �U�    �} t	�E�     �} t	�E�   ��E�    �M�M�}� u&h0hpjj h^  h �j���������u̃}� u3�'���    j h^  h �hh0�r�����   �   �EP�������E��}� u3��   �M�Q���������E��UR�EP�MQj�U�R��������M��U�: u�
���    �
��� �Ej hr  h �hhX�E�P�M�Q�U�P�����P��������} t�M�U��3���]�������������������������������������������������������������������������������������������������������������������������������U���� ��E��=�� u3���   �}� u"�=$� t�����t3���   � ��M��}� ��   �} ��   �UR�#������E��E��8 ��   �M��R������;E���   �E���U����=uo�M�Q�UR�E��Q�U�������uUh�  �U���M��TR�������=�  r&h��hpjj h�   h �j�k�������u̋M���E��D��M����M��O���3���]���������������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E�}� u&hl�hpjj h�   h �j��������u̃}� u3� ���    j h�   h �h��hl��K �����   �%  �U�    �} t�} w�} u�} t	�E�    ��E�   �E��E�}� u&h��hpjj h�   h �j��������u̃}� u3�d���    j h�   h �h��h���������   �   �} t�U� �EP��������E��}� u3��d�M�Q����������U��} u3��F�E�;Mv�"   �5j h�   h �h��h� �U�R�EP�MQ������P�%�����3���]�����������������������������������������������������������������������������������������������������������������U��j�h@�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h��hpjj jNh �j�]�������u̃}� u-����    j jNh �h��h��� �����3���   h�  �UR�]�����=�  s	�E�   ��E�    �E܉E؃}� u#h��hpjj jOh �j�Ӿ������u̃}� u*�(���    j jOh �h��h���v�����3��<j荿�����E�    �UR�������E��E������   �j������ËEԋM�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������U��j�h`�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j蜾�����E�    �EP�MQ�UR�EP�������E��E������   �j������ËE�M�d�    Y_^[��]������������������������������������������������U���EP�MQ�L�����]����������U���EP�MQ�,�����]����������U��Q�E=��  u3��G�M��   }�U���P�M#��&�U�Rj�EPj���u3�f�M��E��U#�]�����������������������������������U���$�} t�} v	�E�   ��E�    �E��E�}� u#hhhpjj jh�j��������u̃}� u0�m���    j jh�hhh�������   �-  �E�    �U�U�} tI�E���t?�U����U��E�;Er�  �M�Uf�f��M���M��:   �E�f��M���M�U�U��}� ��   �E������   �U����U��E�;Er��  �M�U�f�f��M���M�U����U��E����uU����U��E����/t5�U����\t*�M����M��U�;Ur�c  �\   �M�f��U���U�E�E��}� t@�M����t6�E����E��M�;Mr�#  �U�E�f�f�
�U���U�E����E����M�M��}� t�U����t5�M����.t*�E����E��M�;Mr��   �.   �E�f��M���M�U����t6�M����M��U�;Ur�   �E�M�f�f��E���E�M����M����U����U��E�;Ev�e3ɋU�f�
�}�tP�}���tG�E�;Es?�M+M�9h�s�h��U��	�E+E��E�M���Qh�   �U��E�PQ������3���   3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R�C������ _��t3�t	�E�   ��E�    �U��U܃}� u#hP_hpjj jlh�j��������u̃}� u-�B���� "   j jlh�hhP_�������"   ��   ��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���H�E�    �E�    �E�    �} u�e  �} u�} u�} t�} u�H  �} u�} u�} t�} u�+  �} u�}  u�} t�}  u�  �}$ u�}( u�}$ t�}( u��  �}� ��   �E�   �E�E��}� v�M����t�E���E�M����M��܋U����:u2�} t!�}s�  j�MQ�UR�EP�h������M����M�_�} tY3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R�R������E�    �E�    �E�E��	�M����M��U����t4�M����/t�E����\u�U����U���E����.u�U��U�빃}� t>�} t0�E�+E���E��M;M�w�  �U�R�EP�MQ�UR�e������E��E�_�} tY3ɋUf�
�}�tK�}���tB�}v<�E��9h�s�h��M��	�U���U�E���Ph�   �M��Q�R������}� ty�U�;Urq�} t0�E�+E���E��M ;M�w��   �U�R�EP�M Q�UR�������}$ t0�E�+E����E��M(;M�w�   �U�R�E�P�M(Q�U$R�������   �} t0�E�+E���E��M ;M�w�   �U�R�EP�M Q�UR�I������}$ tX3��M$f��}(�tJ�}(���tA�}(v;�U(��9h�s
�h��E��	�M(���M��U���Rh�   �E$��P�?�����3��  �E�   �} t_�} vY3ɋUf�
�}�tK�}���tB�}v<�E��9h�s�h��M��	�U���U܋E���Ph�   �M��Q��������} t_�} vY3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E؋M���Qh�   �U��R�g������} t^�}  vX3��Mf��} �tJ�} ���tA�} v;�U ��9h�s
�h��E��	�M ���MԋU���Rh�   �E��P�������}$ t_�}( vY3ɋU$f�
�}(�tK�}(���tB�}(v<�E(��9h�s�h��M��	�U(���UЋE���Ph�   �M$��Q�������} t	�E�   ��E�    �ỦUȃ}� u&h(hpjj h�   hXj�L�������u̃}� u3�����    j h�   hXh�h(��������   �   �}� t|3�t	�E�   ��E�    �U��U��}� u&h�hpjj h�   hXj�Ǳ������u̃}� u0�����    j h�   hXh�h��g������   ������� "   �"   ��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��=,��t�=,��t�,�P��]��������������U��j j jj jh   @h(�T�,�]�������������U���<�E�    �E�    �E�H��pt	�U��pu'�E�H�U;�u	�E�   ��E�    �E��  �E�H��st�U�B��St	�E�    ��E�   �M��M��U��st�E��St	�E�    ��E�   �M�M��}� u�}� t[�U�;U�uD�E�H�� u	�E�   ��E�    �U�� u	�E�   ��E�    �E�;E�u	�E�   ��E�    �E���  �M�Q��dtv�E�H��itj�U�B��ot^�M�Q��utR�E�H��xtF�U�B��Xt:�M��dt1�U��it(�E��ot�M��ut�U��xt�E��X�,  �M�Q��dtE�E�H��it9�U�B��ot-�M�Q��ut!�E�H��xt�U�B��Xt	�E�    ��E�   �M��dt6�U��it-�E��ot$�M��ut�U��xt�E��Xt	�E�    ��E�   �M�;M�t3��   �U�B%   t	�E�   ��E�    �M��   t	�E�   ��E�    �U�;U�u;�E�H�� t	�E�   ��E�    �U�� t	�E�   ��E�    �E�;E�t3���M�;Uu	�E�   ��E�    �Eċ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE�ǅ ���    ǅ����    ǅ����    ǅ����    ǅ`���    ǅ���    ǅ8���    ǅ����    ǅP���    �EP��h����2���ǅ����    ǅx���    ǅ����    ǅ����    ǅ��������ǅ��������ǅ��������ǅ��������ǅ��������ǅT���    �d����������} tǅ���   �
ǅ���    ����������������� u&h�hpjj h  hx�j觪������u̃����� uI������    j h  hx�h<h��D�����ǅ����������h����t�����������6  �} tǅ����   �
ǅ����    ������������������ u&h��hpjj h  hx�j���������u̃����� uI�P����    j h  hx�h<h��������ǅ���������h��������������16  ǅ����    �U������ǅ����    �����������������������5  ������u������ u��5  ǅ����    ǅd���    ǅT���    ǅ ���    ǅ��������ǅ����    ǅ����    �������Mǅ��������ǅ��������ǅ��������ǅ���������Uf�f������������������U���U����� �N2  ������ �A2  �������� |%��������x��������(����������
ǅ����    ������������k�����	��d�����H�����d�����d�����  �U���%��  �������u\j
��x���Q�UR��������~9��x������$u+������ uh@  j ������R�������ǅ����   �
ǅ����    �������.  j
��x���P�MQ�S���������������x������U������ ��   ������ |#��x������$u������d}ǅ ���   �
ǅ ���    �� ��������������� u&h�hpjj hU  hx�j��������u̃����� uI�]����    j hU  hx�h<h�������ǅ����������h���������������>3  ������;�����~�����������������������������������   ��d�����   3�tǅ����   �
ǅ����    ���������������� u&h��hpjj ha  hx�j��������u̃���� uI�p����    j ha  hx�h<h��������ǅ����������h��������������Q2  ��d����������������I/  �������$�<������� u	������t������u�������u�/  ǅP���   ������Q�UR������P�A  ����.  ǅ���    �������8�����8�����������������`���ǅ����    ǅ��������ǅP���    �.  ������������������ ����������wj�������t��$�\����������������E���������������4���������������#�������ʀ   ����������������������.  ��������*��  ������ u�UR�'������������  j
��x���P�MQ�����������������x������U������ �)  ������ |#��x������$u������d}ǅ���   �
ǅ���    ����������������� u&h �hpjj h�  hx�j薣������u̃����� uI������    j h�  hx�h<h ��3�����ǅ���������h����c����������/  ������;�����~�������� ������������ ����� ����������������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R��������tǅ����   �
ǅ����    ������������������ u&h��hpjj h�  hx�j�7�������u̃����� uI�����    j h�  hx�h<h���������ǅ����������h��������������j.  �v+  �+����������������H�����H���Q藸���������������� }���������������������؉������k�����
�������DЉ������+  ǅ����    ��*  ��������*��  ������ u�UR�������������  j
��x���P�MQ�����������������x������U������ �)  ������ |#��x������$u������d}ǅ����   �
ǅ����    ������������������ u&h��hpjj h�  hx�j臠������u̃����� uI������    j h�  hx�h<h���$�����ǅ����������h����T����������,  ������;�����~��������������������������������������������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R��������tǅ<���   �
ǅ<���    ��<��������������� u&h8�hpjj h�  hx�j�(�������u̃����� uI�z����    j h�  hx�h<h8��������ǅ ���������h���������� ����[+  �g(  �+��������������������������Q舵���������������� }
ǅ���������k�����
�������LЉ������(  ��������(�����(�����I��(�����(���.�D  ��(��������$����E���lu�U���U������   �����������������������   �U���6u,�M�Q��4u �E���E�������� �  �������   �U���3u)�M�Q��2u�E���E������������������e�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu��������   �������ǅd���    �����#�������� ���������������   �������&  ��������0�����0�����A��0�����0���7��#  ��0�������$�̲������%0  u�������� ������ǅP���   ������ u�UR�f�����f��|����   ������ |������d}ǅ����   �
ǅ����    ������������������ u&h��hpjj hz  hx�j��������u̃����� uI�k����    j hz  hx�h<h��������ǅ@���������h���������@����L(  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R�H�������tǅ4���   �
ǅ4���    ��4��������������� u&h��hpjj h~  hx�j��������u̃����� uI�3����    j h~  hx�h<h���~�����ǅ����������h���讴���������'  �w!  �,������������������������Q�A�����f��|����������� ��   ��|���%�   �   k� ��@���ǅ����   ������s������������Ƅ@��� ��h�������P��h���������QtR��@���P������Q��������}
ǅ8���   ��   k� f��|���f������������������ǅ����   �   ������ u�EP�^�������L����  ������ |������d}ǅ����   �
ǅ����    ��������,�����,��� u&h��hpjj h�  hx�j��������u̃�,��� uI�d����    j h�  hx�h<h��������ǅ����������h����߲���������E%  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������P������Qj��������������P�A�������tǅ����   �
ǅ����    ������������������ u&h��hpjj h�  hx�j�ڗ������u̃����� uI�,����    j h�  hx�h<h���w�����ǅ8���������h���觱����8����$  �p  �+��������������������������R�:�������L�����L��� t��L����x u#�p�������������R�F������������d������%   t/��L����Q��������L���� �+���������ǅP���   �(ǅP���    ��L����Q��������L�����������  ��������0  u�������� �������������uǅ����������������������������,��������� u�EP�4������������  ������ |������d}ǅ$���   �
ǅ$���    ��$��������������� u&h��hpjj h:  hx�j��������u̃����� uI�:����    j h:  hx�h<h��������ǅ����������h���赯���������"  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������P������Qj��������������P��������tǅ����   �
ǅ����    ��������|�����|��� u&h��hpjj h>  hx�j谔������u̃�|��� uI�����    j h>  hx�h<h���M�����ǅ����������h����}�����������   �F  �+����������������0�����0���R�������������������� ��   ������ u�p���������������H���ǅ����    ���������������������;�,���}O��H������tB��h��������P��H����R���������t��H�������H�����H�������H�����   ������ u�t�������ǅP���   ��������$�����,�����x�����,�������,�����x��� t��$������t��$�������$���뾋�$���+���������������  ������ u�MQ�©����������  ������ |������d}ǅ���   �
ǅ���    �������t�����t��� u&h��hpjj h�  hx�j�v�������u̃�t��� uI������    j h�  hx�h<h��������ǅ���������h����C���������  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������Q������Rj��������������Q��������tǅ����   �
ǅ����    ��������l�����l��� u&h��hpjj h�  hx�j�>�������u̃�l��� uI�����    j h�  hx�h<h���������ǅp���������h���������p����q  ��  �+����������������(�����(���P螧����������j�������   3�tǅ���   �
ǅ���    �������d�����d��� u&h�hpjj h�  hx�j�X�������u̃�d��� uI�����    j h�  hx�h<h��������ǅh���������h����%�����h����  ��  �������� t�����f������f��������������ǅ8���   �  ǅ���   �������� f��������������@��������������  ������ ��  ������ |������d}ǅ����   �
ǅ����    ��������\�����\��� u&h��hpjj h�  hx�j� �������u̃�\��� uI�r����    j h�  hx�h<h��������ǅ����������h��������������S  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������Q������Rj��������������Q�\�������tǅ���   �
ǅ���    �������T�����T��� u&h(�hpjj h�  hx�j���������u̃�T��� uI�G����    j h�  hx�h<h(�������ǅ`���������h����§����`����(  �  ������������ǅ ���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Yh�  hp�j������]  P��������T�����T��� t ��T�����������������]  �� ����
ǅ�����   ������ u#�E���E�M�Q��A��������������!  ������ |������d}ǅ����   �
ǅ����    ��������L�����L��� u&h��hpjj h  hx�j�H�������u̃�L��� uI�����    j h  hx�h<h���������ǅ ���������h��������� ����{  ������t&h��hpjj h  hx�j�ǋ������u̋������������������������������������Q��A���������������h�������P�����Q������R������P�� ���Q������R������P�   k���0�P��Ѓ���������   t6������ u-��h����4���P������R�   k�	��0�R��Ѓ���������gu;��������   u-��h��������P������R�   ����0�Q��Ѓ����������-u!��������   ��������������������������P萴�����������R  ��������@������ǅD���
   �   ǅD���
   �   ǅ����   ǅ ���   �
ǅ ���'   ǅD���   ��������   t8�   k� �0   f��<����� �����Q�   �� f��<���ǅ`���   �)ǅD���   ��������   t������   �������������� �  �P  ������ u�UR臸�����������������%  ������ |������d}ǅ����   �
ǅ����    ��������D�����D��� u&h��hpjj h�  hx�j��������u̃�D��� uI�T����    j h�  hx�h<h��������ǅX���������h����Ϣ����X����5  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R�1�������tǅ����   �
ǅ����    ������������������ u&h�hpjj h�  hx�j�ʇ������u̃����� uI�����    j h�  hx�h<h��g�����ǅ���������h���藡���������  �`  �1����������������P�����P���Q�]�������������������  ��������   �P  ������ u�EP�%������������������%  ������ |������d}ǅ����   �
ǅ����    ������������������ u&h��hpjj h�  hx�j蠆������u̃����� uI������    j h�  hx�h<h���=�����ǅ���������h����m����������  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������P������Qj��������������P�ϸ������tǅ����   �
ǅ����    ������������������ u&h��hpjj h�  hx�j�h�������u̃����� uI�����    j h�  hx�h<h��������ǅ����������h����5����������  ��  �1��������������������������R��������������������z	  �������� ��  ��������@�T  ������ u�UR脛�������������������'  ������ |������d}ǅ����   �
ǅ����    ������������������ u&h��hpjj h�  hx�j�0�������u̃����� uI�����    j h�  hx�h<h���������ǅ����������h���������������c  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R�_�������tǅ����   �
ǅ����    ������������������ u&h��hpjj h�  hx�j���������u̃����� uI�J����    j h�  hx�h<h��������ǅ����������h����Ŝ���������+  �	  �3��������������������������Q�X��������������������S  ������ u!�UR�0���������������������)  ������ |������d}ǅx���   �
ǅx���    ��x�����p�����p��� u&h��hpjj h�  hx�j�ځ������u̃�p��� uI�,����    j h�  hx�h<h���w�����ǅ����������h���觛���������  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R�	�������tǅh���   �
ǅh���    ��h�����`�����`��� u&h��hpjj h  hx�j袀������u̃�`��� uI������    j h  hx�h<h���?�����ǅ����������h����o�����������  �8  �5����������������|�����|���Q����������������������  ��������@�R  ������ u�EP�ɖ������������������&  ������ |������d}ǅX���   �
ǅX���    ��X�����P�����P��� u&h��hpjj h  hx�j�v������u̃�P��� uI������    j h  hx�h<h��������ǅt���������h����C�����t����  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������P������Qj��������������P襱������tǅH���   �
ǅH���    ��H�����@�����@��� u&h��hpjj h  hx�j�>~������u̃�@��� uI�����    j h  hx�h<h���ۼ����ǅl���������h���������l����q
  ��  �2����������������d�����d���R螔������������������O  ������ u�EP�w�����3ɉ������������'  ������ |������d}ǅ8���   �
ǅ8���    ��8�����0�����0��� u&h��hpjj h4  hx�j�#}������u̃�0��� uI�u����    j h4  hx�h<h���������ǅ\���������h���������\����V	  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������Q������Rj��������������Q�R�������tǅ(���   �
ǅ(���    ��(��������������� u&h��hpjj h8  hx�j��{������u̃����� uI�=����    j h8  hx�h<h��舺����ǅT���������h���踕����T����  �  �3����������������L�����L���P�K�����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�X�����\�����������   ���������������X�����������\����������� �  u(������%   u��X�����\����� ��X�����\��������� }ǅ����   �%���������������������   ~
ǅ����   ��X����\���u
ǅ`���    �   i��  ��������������������D�������������������D��� ��X����\�����   ��D����RP��\���R��X���P蚓����0��4�����D����RP��\���Q��X���R�֑����X�����\�����4���9~��4���� �����4�����������4�������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0��������������������u������ u�  ��8��� �a  ��������@��   ��������   t!�   k� �-   f��<���ǅ`���   �V��������t!�   k� �+   f��<���ǅ`���   �*��������t�   k� �    f��<���ǅ`���   ������+�����+�`�����������������u������Q�UR������Pj ��  ��������Q������R�EP��`���Q��<���R��  ����������t'��������u������R�EP������Qj0�l  ����P��� ��   ������ ��   �����������������������������<�����������������<��� ��   ��h����z���P��h����n���� �HtQ�����R��|���P�r����������������� ǅ���������2������Q�UR��|���P�)  ������������������X����(������R������P�MQ������R������P�  �������� |'��������t������R�EP������Qj �8  ����T��� tj��T���R������ǅT���    ������d��� t��d���tǅ����    �
ǅ����   ������������������ u&hh�hpjj h�  hx�j�v������u̃����� uI�T����    j h�  hx�h<hh�蟴����ǅ4���������h����Ϗ����4����5  �������  ������ ��  ǅ����    ���������������������;�������  ��������������������������������������   ������$�@����������E�������MQ�������d  ���������E�������MQ�ŋ�����@  ���������E�������MQ�ԣ�����  ���������E�������MQ谣������   ���������E�������MQ�Y�������   ���������E�������MQ�k������������������   3�tǅ����   �
ǅ����    ������������������ u&h��hpjj h2	  hx�j��s������u̃����� uF�C����    j h2	  hx�h<h��莲����ǅ,���������h���辍����,����'����������������$�����h���蕍����$����M�3��5�����]��V���;�;�J�7��������'�6� �I ����t����� ����{�����D����q��b�����   	
���ǰ��c�3�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E�H��@t�U�z u�E����U�
�4�EP�MQ�������Ё���  u�E� ������M����E�]�������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�U������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��~�U�    �E�E��M���M�}� ~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������뛋E�8 u�M�U���]����������������������������������������������U���  ���3ŉE�ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    �EP��d����rk��ǅ����    �������P����} tǅ0���   �
ǅ0���    ��0�����`�����`��� u&h�hpjj h  hx�j�Aa������u̃�`��� uI蓧���    j h  hx�h\h��ޟ����ǅ���������d����{��������  �} tǅ(���   �
ǅ(���    ��(����� ����� ��� u&h��hpjj h  hx�j�`������u̃� ��� uI�����    j h  hx�h\h���5�����ǅ���������d����ez���������  ǅ����    ǅ����    ǅ����    ǅ����    ǅt���    �Uf�f������������������U���U����� ��  ������ ��  �������� |%��������x��������(�����<����
ǅ<���    ��<���������k�����	��������H�����������������   3�tǅ8���   �
ǅ8���    ��8�����T�����T��� u&h��hpjj he  hx�j�_������u̃�T��� uI�b����    j he  hx�h\h��譝����ǅ����������d�����x���������n  ��������,�����,�����  ��,����$�h�ǅ����   ������Q�UR������P�  ���J  ǅ����    ������������������������������������ǅ����    ǅ��������ǅ����    ��  �������������������� ������������wj�����������$������������������E���������������4���������������#�������ʀ   ����������������������e  ��������*u:�UR�Ot���������������� }���������������������ى������k�����
�������LЉ������  ǅ����    ��  ��������*u'�EP��s���������������� }
ǅ���������k�����
�������DЉ������  ��������������������I������������.�1  �����������$����U���lu�M���M��������   �����������������������   �M���6u+�E�H��4u�U���U������ �  �������   �M���3u(�E�H��2u�U���U������%����������S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    ������#�������� ���������������   �������D  ��������������������A������������7��
  ��������4��$�����������0  u�������� ������ǅ����   �EP��q����f�������������� ��   ���������   �   k� ������ǅL���   ��L���s��}�����L���Ƅ���� ��d���谧��P��d���褧��� �HtQ������R������P訞������}
ǅ����   ��   k� f������f������������������ǅ����   �s	  �UR��p���������������� t�������x u#�p�������������R�������������d������%   t/�������Q������������� �+���������ǅ����   �(ǅ����    �������Q���������������������  ��������0  u�������� �������������uǅ4���������������4�����4����������EP��o������������������ ��   ������ u�p�������������������ǅ����    ���������������������;�����}O���������tB��d����ƥ��P�������P�Ӧ������t������������������������������   ������ u�t�������ǅ����   ������������������������������������������ t���������t��������������뾋�����+��������������2  �UR�n������\���膏������   3�tǅD���   �
ǅD���    ��D�����$�����$��� u&h�hpjj h�  hx�j�tW������u̃�$��� uI�Ɲ���    j h�  hx�h\h�������ǅ ���������d����Aq���� �����	  �g  �������� t��\���f������f����\����������ǅ����   �-  ǅ����   �������� f��������������@������������������ǅt���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Yh�  hp�j������]  P�3R���������������� t ��������������������]  ��t����
ǅ�����   �E���E�M�Q��A���������������d�������P������Q������R������P��t���Q������R������P�   k���0�P��Ѓ���������   t6������ u-��d����~���P������R�   k�	��0�R��Ѓ���������gu;��������   u-��d����7���P������R�   ����0�Q��Ѓ����������-u!��������   ��������������������������P��~������������  ��������@������ǅ����
   �   ǅ����
   �   ǅ����   ǅ����   �
ǅ����'   ǅ����   ��������   t8�   k� �0   f��������������Q�   �� f������ǅ����   �)ǅ����   ��������   t������   �������������� �  t�UR�ނ�����������������   ������%   t�MQ贂�����������������   �������� tE��������@t�MQ�Nj��������������������UR�2j��������������������@��������@t�MQ�	j�������������������UR��i����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ������������������ }ǅ����   �%���������������������   ~
ǅ����   �����������u
ǅ����    �   i��  ������������������������������������������ �������������   �������RP������R������P�=k����0�������������RP������Q������R�yi��������������������9~���������������������������������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0�������������������� �a  ��������@��   ��������   t!�   k� �-   f������ǅ����   �V��������t!�   k� �+   f������ǅ����   �*��������t�   k� �    f������ǅ����   ������+�����+�������x�����������u������Q�UR��x���Pj �	  ����P���Q������R�EP������Q������R��	  ����������t'��������u������R�EP��x���Qj0�F	  �������� ��   ������ ��   ��������|����������������������������������������������� ��   ��d����4���P��d����(���� �HtQ��|���R������P�,�������X�����X��� ǅ���������2������Q�UR������P�  ����|����X�����|����X����(��P���R������P�MQ������R������P�  �������� |'��������t������R�EP��x���Qj �  �������� tj������R��\����ǅ����    ���������� t������tǅH���    �
ǅH���   ��H�����@�����@��� u&hh�hpjj h�  hx�j�M������u̃�@��� uF�����    j h�  hx�h\hh��Y�����ǅ���������d����g���������������������d����jg��������M�3��
l����]Ð�;��� �������A����������� �I [���*�<� ���~�3�1�������������'�P��=���   	
��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E�H��@t�U�z u�E����U�
�4�EP�MQ�������Ё���  u�E� ������M����E�]�������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�U������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��~�U�    �E�E��M���M�}� ~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������뛋E�8 u�M�U���]����������������������������������������������U���4���3ŉE�V�E�H��@�d  �UR�?x�������t@�EP�.x�������t/�MQ�x���������UR�x���������P��E���E���E��H$�����у�tj�EP��w�������t@�MQ��w�������t/�UR�w���������EP�w���������P��E���E���MԊQ$������uh�M�Q���U�E�M�H�}� |2�U�f�Mf��U����  f�U�E����U�
f�E��  ��EP�MQ�h�����  �(  �UR�w�������t@�EP��v�������t/�MQ��v���������UR��v���������P��E���E���E��H��   ��   �URj�E�P�M�Q迊������t
���  ��   �E�    �	�U����U��E�;E�}s�M�Q���U؋E�M؉H�}� |.�U��M��T��E�����   �U�E����U�
��EP�M��T�R�������E�}��u���  �k�|����E%��  �[�E�H���M܋U�E܉B�}� |/�M�f�Ef��M����  f�M�U����M�f�E����UR�EP�f����^�M�3���`����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    3�f�E�} t	�E�   ��E�    �M܉M؃}� u#h��hpjj j3h�j��@������u̃}� u-�3����    j j3h�h�h����������  �M�E�E��M�Q��v�����E�    �U�R�EP������f�E��E������   ��M�Q�}�����f�E�M�d�    Y_^[��]��������������������������������������������������������������������U��EP�MQ�e����]�����������U����E�E�M�M��E�    �	�U����U��}�}�E��M���E����E��M���M��Ӌ�]���������������������U��Q�E�    �	�E����E��}�}�M��U��    ���]������������������U����E�������E��E%  �yH���@�   +ȉM��   �M���U��E��M��R�E�P�M��U��P�RH�����E��M����M��	�U����U��}� |)�}� t#�E��M��Rj�E��M��R�H�����E��ȋE���]���������������������������������������������������������U��Q�E�    �	�E����E��}�}�M��U�<� t3���߸   ��]��������������������������U����E�    �E���E��M����M�E��������E��U��  �yJ���B�   +E�   �M���U�E��M��#U�t'�E�P�MQ�k������u�U�R�EP�<j�����E����M���E��M#��E��M���U����U��	�E����E��}�}�M��U��    ��E��]�������������������������������������������������������������U���V�E�������E��E%  �yH���@�E�����M����҉U��E�    �E�    �	�E����E��}�}M�M��U��#E�E�M��U���M���M��U���E��M��U�E��M���    +M��U���U���E�   �	�E����E��}� |.�M�;M�|�U�+U��E��M�u������E��M��    ��^��]���������������������������������������������������������������������U����E�������E��E%  �yH���@�   +ȉM�����M����҉U�E��M��#U�t3��1�E����E��	�M����M��}�}�U��E�<� t3���߸   ��]�����������������������������������������������U����E�    �EE�E��M�;Mr�U�;Us	�E����E��M�U���E���]�������������������U���@���3ŉE��E�H
���  ���?  �M��U�B
% �  �E��   k� �E�H�L�   �� �E�H�L��U����   ��D��}����u8�E�    �U�R�{T������t	�E�    ��E�P�X�����E�   �  �M�Q�U�R�������E��E̋M�QR�E�P��s������t	�M����M��U�E�J+H9M�}�U�R�W�����E�    �E�   �  �E�M�;Hn�U�R�E�P�z������M̉M��U�B+E��EȋM�Q�U�R��u�����E�HQ�U�R�ls�����E�H��Q�U�R��u�����E�    �E�   �   �E�M�;|T�U�R�W�����   k� �T���   ��   k� �T��U�BP�M�Q�mu�����U��MA�E��E�   �C�U�E�B�Eع   k� �D�%����   k� �D��E�HQ�U�R�u�����E�    �E�H���    +щUă}� t	�E�   ���E�    �   k� �E؋M���D�EԉEЋM�y@u�U�EЉB�   �� �U�D����M�y u�U�EЉ�E܋M�3���V����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��h0��EP�MQ�~����]�������U��hH��EP�MQ�u~����]�������U������3ŉE��E�    �E�H
���  f�M�U�B
% �  f�E�   k� �E�H�L�   �� �E�H�L��U����   ��D�j@�U�R�p������t�   k� �D�   �f�U�f��f�U��E�=�  u�E�   �   k� �E�L��H�   �� �E�L���U��E�ЋMf�Q�E�M�3���T����]����������������������������������������������������������������������������U������3ŉE��EPj j j �MQ�UR�EP�M�Q��s���� �E�UR�E�P��n�����E�}�u	�M���M�E�M�3��IT����]�����������������������������������������U���T���3ŉE�3�f�E��E�    �E�    �E�    �E�    �Mf�Q
f�U�Ef�H
f�M��U��E�3Ё� �  f�U��M���  f�M��U���  f�U��E��M��f�E��U���  }�E�=�  }�M����  ~9�U���t	�E� �����E� ���E�M��H�U�B    �E�     �  �M���?  "�U�B    �E�@    �M�    ��  �U��u9f�E�f��f�E�M�Q�����u�E�x u�M�9 u3ҋEf�P
�  �M��uMf�U�f��f�U�E�H�����u3�U�z u*�E�8 u"�M�A    �U�B    �E�     �R  �E�    �E�    �	�M؃��M؃}���   �U���U��E�   �   +E؉E��	�Mȃ��Mȃ}� ~x�UỦU��EEԉE��M܍T��U��E���U���ȉM��M�Q�U�R�E��Q�<�����E��}� t�U�f�D�f���M�f�D�Ũ��ŰEԃ��E��y����M܃��M��<����U���?  f�U��E��~%�M���   �u�U�R�(9����f�E�f��f�E����M��Qf�U�f��f�U��E��},�M���t	�UЃ��UЍE�P��1����f�M�f��f�M��̃}� t�U���f�U��E�= �  �M����� �� � u_�}��uP�E�    �}��u8�E�    �U�����  u� �  f�E�f�M�f��f�M��f�U�f��f�U��	�E����E��	�M���M��U���  |6�E���t	�E� �����E� ���M�UĉQ�E�@    �M�    �-�Uf�E�f��M�U�Q�E�M��H�U��E�ЋMf�Q
�M�3��P����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U������3ŉE��p���`�E�} u�   �} }�M�ىM�����`�U�} u3��Mf��} tp�U��T�U�E���E�M���M�}� u��kU�U�U�E���� �  |#�U��E��J�M�R�U��E���E�M��M�U�R�EP�rq����늋M�3��@N����]����������������������������������������������������������������U����E���   �t	�E�   ��E�    �U��U�E�H��   �t	�E�   ��E�    �U��U��E���U�
�E�H��M�U�J�E�H��M��U�J��]����������������������������������U����E�H��t	�E�   ���E�    �U��U�E�H��t	�E�   ���E�    �U��U��E�H��U�J�E�H��M�U�J�E���M��U�
��]���������������������������������������U���   ���3ŉE��E��E�3�f�M�ǅl���   �E�    �E�    �E�    ǅp���    �E�    ǅ|���    �E�    �E�    �E�    �E�    3�f�U�3�f�E��E�    �E�    �}$ tǅh���   �
ǅh���    ��h�����\�����\��� u#h�hpjj j~hj�-������u̃�\��� u-�hs���    j j~hh�h��k����3��  �E�E̋M̉M��	�Ũ��ŰE���� t!�U����	t�M����
t�E����u�Ƀ}�
�;  �Ů�EӋM̃��M̋Uȉ�`�����`����  ��`����$���MӃ�1|�UӃ�9�E�   �Ẽ��E��   �MӋU$����   ��;�u	�E�   �`�Eӈ�t�����t���+t��t���-t#��t���0t�*�E�   �1�E�   3�f�M��"�E�   � �  f�U���E�
   �Ẽ��E��U  �E�   �MӃ�1|�UӃ�9�E�   �Ẽ��E��|�MӋU$����   ��;�u	�E�   �[�EӉE��M���+�M��}�:w5�U�����$���E�   �+�E�   �"�M̃��M��E�   ��E�
   �Ũ��U��  �EӃ�1|�MӃ�9�E�   �Ũ��U��K�EӋM$����   ��
;�u	�E�   �*�Uӈ�T�����T���0t�	�E�   ��E�
   �E��E��5  �E�   ��M̊�UӋẼ��E��MӃ�0|:�UӃ�91�}�s �E����E��MӃ�0�U��
�E����E��	�M����M���UӋE$����   ��;�u	�E�   �R�MӉM��U���+�U��}�:w,�E����$��E�   �"�Ũ��U��E�   ��E�
   �Ẽ��E��`  �E�   �E�   �}� u'��M̊�UӋẼ��E��MӃ�0u�U����U�����E̊�MӋŨ��U��EӃ�0|8�MӃ�9/�}�s'�U����U��EӃ�0�M���U����U��E����E���MӉM��U���+�U��}�:w,�E���X�$�L�E�   �"�Ũ��U��E�   ��E�
   �Ẽ��E��z  �E�   �MӃ�0|�UӃ�9�E�   �Ẽ��E���E�
   �M��M��=  �Ũ��U��EӃ�1|�MӃ�9�E�	   �Ũ��U��X�Eӈ�x�����x���+t0��x���-t��x���0t�%�E�   �)�E�   ǅl���������E�   ��E�
   �M��M��  ǅp���   ��Ů�EӋM̃��M��UӃ�0u���EӃ�1|�MӃ�9�E�	   �Ũ��U���E�
   �Ẽ��E��R  �MӃ�1|�UӃ�9�E�	   �Ẽ��E��*�Mӈ�X�����X���0t�	�E�   ��E�
   �U��U���   ǅp���   �E�    ��E̊�MӋŨ��U��EӃ�0|,�MӃ�9#kU�
�EӍLЉM��}�P  ~	�E�Q  �뺋U��U���E̊�MӋŨ��U��EӃ�0|�MӃ�9���E�
   �Ũ��U��g�}  tQ�Ẽ��E��Mӈ�d�����d���+t��d���-t��E�   ǅl���������E�   ��E�
   �U��U���E�
   �Ẽ��E������M�Ủ�}� �`  �}� �V  ��|��� �I  �}�vF�   k��T���|�   k��T����   k��T��E�   �U����U��E����E��}� ��   �M����M��	�U����U��E����u�U����U��E����E��ٍM�Q�U�R�E�P�T������l��� }�M��ىM��U�U��U���p��� u	�E�E�E��}� u	�M�+M�M��}�P  ~	�E�   �E�}�����}ǅ|���   �0�UR�E�P�M�Q�vZ����f�U�f�U��E։E��MډM�f�U�f�U��3�f�E�3�f�M��UĉU��E��E��}� u$3�f�M�3�f�U��EĉE��M��M��U����U��Y�}� t(��  f�E��E�   ��E�    3�f�M��U����U��+��|��� t"3�f�E�3�f�M��UĉU��E��E��M����M��Uf�E�f��M�U��Q�E�M��H�U��E�ЋMf�Q
�E��M�3���B����]Ë�L���������������O�N���~�l�u���  �������  �������  �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE��M  f�E��M   f�M���   f�U��E��C�E���E���E���E���E���E���E���E���E���E���E���E�?�E�   f�Ef�EЋM�M��U�U��E�% �  f�E��MЁ��  f�M��U̅�t	�E�@-��M�A �UЅ�uj�}� ud�}� u^3��Mf��Ú� �  u	�E�-   ��E�    �E�M��H�U�B�   k� �U�D
0�   �� �M�D �   ��  �UЁ��  �b  �   �Mf��}�   �u�}� tP�U���   @uEj jvh�hh0h�j�E��P�of����P�)�����M�A�E�    ��   �U̅�tT�}�   �uK�}� uEj j|h�hh�h�j�E��P�f����P�G)�����M�A�E�    �   �}�   �uK�}� uEj h�   h�hh�hDj�U��R�e����P��(�����E�@�E�    �Cj h�   h�hhPh�j�M��Q�we����P�(�����U�B�E�    �\  �E���f�E��MЁ��   f��|����U���f�U��E��M����U��M�����U��M����+E��E��U���f�U�f�E�f�E��M��M��U��U�3�f�E�j�M���Q�U�R�R�����E�=�?  |f�M�f��f�MȍU�R�E�P��^�����Mf�U�f��E��tn�M�M�M�} ^3ҋEf��Ḿ� �  u	�E�-   ��E�    �U�E��B�M�A�   k� �M�D0�   �� �E�D �   �.  �}~�E   �M����?  �M�3�f�U��E�    �	�E����E��}�}�M�Q��"������}� }-�U��ځ��   �U��	�E����E��}� ~�M�Q�y������U���UԋE���E��	�M����M��}� ~a�U��U؋E�E܋M��M��U�R�M"�����E�P�A"�����M�Q�U�R������E�P�%"�����M���0�UԈ
�Eԃ��E��E� 됋Mԃ��MԋUԊ�EǋMԃ��M��Uǃ�5|_�	�Eԃ��EԋM��9M�r�U����9u�M��0�ًU��9U�s�Eԃ��EԋMf�f���Ef��MԊ���EԈ�   �	�Mԃ��MԋU��9U�r�E����0u�ߋU��9U�s[3��Mf��Ú� �  u	�E�-   ��E�    �E�M��H�U�B�   k� �U�D
0�   �� �M�D �   �&�U���E�+��M�A�U�B�M�D �E��M�3��9����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EP�M�R�E�Q�"�����E��}� t0�U��Rj�E�HQ��!�����E��}� t�U�B���M�A�U��R�E�HQ�U�BP�!�����E�}� t�M�Q���E�P�M��Q�U�BP�M�QR�!������]����������������������������������������������������U����E�    �E%�   t	�M����M��U��   t	�E����E��M��   t	�U����U��E%   t	�M����M��U��   t	�E����E��M��   t�U���   �U��E% `  �E��}� @  w�}� @  t$�}� t�}�    t#�:�}� `  t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��@�  �U�}�@t!�}� �  t&�}�@�  t�'�E�   �E���M���   �M���U���   �U��E���]�����������������������������������������������������������������������������������������������U��Q�E�    �E��?th�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]�����������������������������������������������U��Q�]��e���U��E�P�7�������]�����������������U����} t^��}��E�P�F  ���E��M#M�U��#U�ʉM�E�;E�t'�M�Q�,  ��f�E��m���}��U�R�  ���E�E�M��} t)�=@�|�UR�EP�J   ���M��	�U�    �   ��]�����������������������������������������������U����E%�E�]��M�Q�������E��U#U�E��#E�ЉU�M�;M�u�E��+�U�R�s   ���E��E�P�g�����]��M�Q�D�������]������������������������������U��Q�E��  �E�P�������]����������������������U����E�    �E��t�M��ɀ   �M��U��t�E�   �E��M��t�U���   �U��E��t�M���   �M��U��t�E�   �E��M��   t�U���   �U��E%   �E��}�   w�}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U��� @  �U���E�    �E���M��� `  �M��U��   �U�}�   t�}�   t�}�   t�$�E�@�  �E���M���@�M���U��� �  �U��E���]�����������������������������������������������������������������������������������������������U��Q�s9���E��E�P���������]���������������������U����E�    �E��t	�M����M��U��t	�E����E��M��t	�U����U��E��t	�M����M��U�� t	�E����E��M��t�U���   �U��E%   �E��}�   �}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��   �U�t*�}�   t�}�   t�"�E��E���M���   �M���U���   �U��E%   t�M���   �M��E���]�����������������������������������������������������������������������������������������U��Q�E�    �E��?tn�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]����������������������������������������U��QV�}���=@�|�E�P�3����������������M�Q������^��]������������������U�����}��E�P�L������E�M#M�U��#U�ʉM�E�;E�t'�M�Q�2  ��f�E��m���}��U�R�
������E�=@�|B�EP�MQ�^������E��U�#��E�#�;�t�E�E�   ����E�E����E��]���������������������������������������������������U��E%����P�MQ��3����]�������U����7��� �E����jV���D����}� t/�M��Q�%  t �M��Q���U��E��@    �M��A��  ��]����������������������������U���3�f�E��M��t�U���f�U��E��t�M���f�M��U��t�E���f�E��M��t�U���f�U��E��t�M��� f�M��U��   t�E���f�E��M��   �M��}�   w�}�   t&�}� t�}�   t&�B�}�   t+�7f�U�f�U��-�E�   f�E���M���   f�M���U���   f�U��E%   �E�t�}�   t�}�   t"�(�M���   f�M���U���   f�U��f�E�f�E��M��   t�U���   f�U�f�E���]�����������������������������������������������������������������������������������������������������U����} 	 u>�}�u8��}��E�%=  ==  u$�=@�|�]��M�����  ���  u�;��7j hN  h�hh@�U������R�EPj �����P�������]�����������������������������������������U�����}��E�P�������E��=@�|�]�M�Q������E���E���]������������������U��Q�} t��}��E�P�������M��} t
������U���]�����������������������������U��EP�����]����������������U��j
j �EP�Q2����]������������U��EPj
j �MQ������]��������U��EP�MQ�<>����]������������U��j
j �EP�6����]������������U��EPj
j �MQ�;����]��������U��j
j �EP�1����]������������U��EPj
j �MQ�I����]��������S�܃������U�k�l$���@�=@�}M�C���t�S��K;�t�S���S�݋C��S;�u�C�E���E�    �E��  ��   �Kfn�fE��pE� fE�fpE� fEЋS���  ���  ��   �C�o fE�foE�f�E�fE�foE�fuE�fE�foE�fuE�fE�foE�f�E�fE�foE�f�ȉM��}� t2�U��U��E�C�C�K��C;�u�K�M���E�    �E��:�S���S�*�C��S;�u�C��C���u3���S���S�%�����]��[�������������������������������������������������������������������������������������������������������������SV�L$�T$�\$������tQ+���   t�
:uH��D�B��v4��u�
%�  =�  wً
;u҃�v����������#Ʃ����t�3�^[Íd$ ���^[�����������������������������������������U����=4� ��  �} t	�E�   ��E�    �E��E��}� u&hԸhpjj h�   h�j�������u̃}� u3�cM���    j h�   h�hthԸ�E���������0  �} t	�E�   ��E�    �U�U��}� u&hp�hpjj h�   h�j�������u̃}� u3��L���    j h�   h�hthp��-E���������   �}���w	�E�   ��E�    �M�M�}� u&hLhpjj h�   h�j�	������u̃}� u0�^L���    j h�   h�hthL�D���������.�EP�MQ�UR�������j �EP�MQ�UR�N������]�������������������������������������������������������������������������������������������������������������������������U���L�} �n  �EP�M������} t	�E�   ��E�    �M��M�}� u#hԸhpjj j;h�j��������u̃}� u=�K���    j j;h�h0hԸ�kC�����E�����M�����E���  �} t	�E�   ��E�    �E��E�}� u#hp�hpjj j<h�j�@������u̃}� u=�J���    j j<h�h0hp���B�����E�����M�����E��T  �}���w	�E�   ��E�    �U�U�}� u#hLhpjj j=h�j�������u̃}� u=�
J���    j j=h�h0hL�XB�����E�����M�����E���   �M��P����   �⃼�    u)�EP�MQ�UR�������EЍM��L���E��   �m�E��M̍M��:P��P�U�R�,�����E��E���E�M��UȍM��P��P�E�P��+�����E��M���M�U���Ut�}� t�E�;E�t��M�+M��MčM������E��3���]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�RP�EP�������E��}� u	�E�    ��E������E���]�������������������������U���DV�E�    �E�    �E�    jj j �EP�(�����EĉUȋM�#Mȃ��t#jj j �UR�(�����ẺUЋE�#EЃ��u�G��� �2  �M+M̋UUЉM܉U��}� �?  
�}� �3  h   j�(P�$�E��}� u%�QG���    �E�   �E������E�������   h �  �EP�/"�����E�}� |	�}�   r	�E�   ��M܉M��U��U��}� |	�}�   r	�E�   ��E܉E�M�Q�U�R�EP� ������E��}��u(����8u�F���    �E�   �E���EԉU��*�E���M�+ȋE�M܉E��}� �W���|
�}� �K����M�Q�UR�g!�����E�Pj �(P��   �}� ��   |
�}� ��   j �MQ�UR�EP��&�����EԉU؋M�#M؃��t]�UR�s	����P�X��t	�E�    ��E������E虉EԉU؋E�#E؃��u!��E���    �E�   ��������0�M�#M؃��t'j �U�R�E�P�MQ�W&�����E��U��U�#U����u	�oE��� �3�^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u�^���     �	   �b  �} |�E;\�s	�E�   ��E�    �M��M܃}� u#hhbhpjj j7h�j��������u̃}� u;�����     �D��� 	   j j7h�h�hhb�O<�����	   ��  �E���M������P��D
��t	�E�   ��E�    �M؉Mԃ}� u#hdchpjj j8h�j��������u̃}� u;�S���     �aC��� 	   j j8h�h�hdc�;�����	   �1  �} |�} r	�E�   ��E�    �EЉẼ}� u#h	hpjj j9h�j��������u̃}� u;�����     ��B���    j j9h�h�h	�!;�����   �   �UR�|G�����E�    �E���M������P��D
��t�MQ�UR�EP�1�����E��93�u#h(ahpjj jAh�j���������u��0B��� 	   �E�	   �E������   ��EP�Z�����ËE�M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u&hphpjj h�   h8
j��������u̃}� u0��@���    j h�   h8
h�hp�+9�����   ��U�,��3���]���������������������������������������������U����} @  t�} �  t�}   t	�E�    ��E�   �E��E��}� u&h�
hpjj h�   h8
j��������u̃}� u0�@���    j h�   h8
hTh�
�V8�����   ��U�,��3���]��������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} @  t-�} �  t$�}   t�}   t�}   t	�E�    ��E�   �E��E܃}� u#h(	hpjj j6h8
j��������u̃}� u.��>���    j j6h8
h�
h(	�97���������  �}�u�>��� 	   ����  �} |�U;\�s	�E�   ��E�    �E؉Eԃ}� u#h`hpjj j9h8
j���������u̃}� u.�N>��� 	   j j9h8
h�
h`�6��������2  �U���E������P��T��t	�E�   ��E�    �EЉẼ}� u#h�`hpjj j:h8
j�f�������u̃}� u.�=��� 	   j j:h8
h�
h�`�	6��������   �UR�fB�����E�    �E���M������P��D
��t�MQ�UR�^�����E��9�E=��� 	   3�u#h(ahpjj jEh8
j��������u��E������E������   ��UR�H�����ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E���M������P��D
%�   �E��M���U������P��L$�����щU�E�E��}�   $�}�   �a  �}� @  tm�}� �  t$�  �}�   �=  �}�   ��   �  �M���U������P��L������U���E������P��L�`  �E���M������P��D
�   �M���U������P��D�U���E������P��T$�​E���M������P��T$��   �M���U������P��L�ɀ   �U���E������P��L�E���M������P��D
$$��M���U������P��D$�u�U���E������P��T�ʀ   �E���M������P��T�M���U������P��L$�က��U���E������P��L$�}� u� �  ��}� u	� @  ���   ��]�������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��L���3�P�E�d�    �EP�M��]����E�    �} t�M�U��} t	�E�   ��E�    �E��E܃}� u#h�hpjj j^h�j�>�������u̃}� uD�8���    j j^h�h<h���0�����E�    �E������M�����E��  �} t�}|�}$~	�E�    ��E�   �U؉Uԃ}� u#hPhpjj j_h�j��������u̃}� uD��7���    j j_h�h<hP�F0�����E�    �E������M��u���E��s  �M�M��E�    �U��E�M���M�M��P>����t-�M��D>����zt~�M��4>��Pj�E�P������E��j�M�Q�M��>��P�������EЃ}� t�U��E�M���M���U��-u�E���E�M��U�E���E���M��+u�U��E�M���M�} |�}t�}$~.�} t�U�E��E�    �E������M��m
���E��k  �>�} u8�M��0t	�E
   �&�U����xt�M����Xu	�E   ��E   �} u8�E��0t	�E
   �&�M����xt�E����Xu	�E   ��E   �}u9�U��0u0�E����xt�U����Xu�M���M�U��E�M���M�����3��u�E�j�U�R�M��<��P�@�������t�E��0�E��Qh  �M�Q�M��j<��P��������t0�U��a|�E��z�M�� �M���U�ŰẼ�7�E���f�M�;Mr�\�U���U�E�;E�r�M�;M�u���3��u9U�w�U��UU�U���E���E�} u��M��U�E���E��!����M���M�U��u�} t�E�E��E�    �f�M��u*�U��uV�E��t	�}�   �w�M��u=�}����v4�4��� "   �U��t	�E�������E��t	�E�   ���E�����} t�M�U��E��t�M��ىM�U�U��E������M������E��M�d�    Y��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�EP������]������������������U��j�EP�MQ�UR�EP������]������������������U��=4� uj �EP�MQ�URh��L�������j �EP�MQ�URj �0�����]����������������������������U��=4� uj�EP�MQ�URh����������j�EP�MQ�URj �������]����������������������������U��EP�MQ�URh�]�����]�������������������U��EPj �MQhsa�[����]���������������������U��EP�MQ�URhsa�)����]�������������������U��EP�MQ�URh``������]�������������������U��EPj �MQh�]������]���������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �1"���    �� ��E��E�    �} t	�E�   ��E�    �U��U܃}� u#h��hpjj j4h�j���������u̃}� u+�P0���    j j4h�hh���(��������i�M�Q� �����E�    �U�R������EԋEP�MQ�UR�E�P�U���E؋M�Q�U�R�,�����E������   ��E�P�&����ËE؋M�d�    Y_^[��]���������������������������������������������������������������������������������������U��EPj �MQh``�����]���������������������U��j�h�d�    P��lVW���3�P�E�d�    �EP�M��[����E�    �} t�M�U��} t	�E�   ��E�    �E�E��}� u#h�hpjj jch@j�<�������u̃}� uN�.���    j jch@h�h���&�����E�    �E�    �E������M�����E��U��<  �} t�}|�}$~	�E�    ��E�   �U܉U؃}� u#hPhpjj jdh@j��������u̃}� uN��-���    j jdh@h�hP�:&�����E�    �E�    �E������M��b���E��U��  �M�M��E�    �E�    �U��E�M���M�M��34����t-�M��'4����zt~�M��4��Pj�E�P�������E��j�M�Q�M���3��P�������Eԃ}� t�U��E�M���M���U��-u�E���E�M��U�E���E���M��+u�U��E�M���M�} u8�U��0t	�E
   �&�E����xt�U����Xu	�E   ��E   �}u9�M��0u0�U����xt�M����Xu�E���E�M��U�E���E�E�RPj�j�������E��U�j�M�Q�M���2��P��������t�U��0�U��Th  �E�P�M���2��P�n�������t0�M��a|�U��z�E�� �E���M�MЋUЃ�7�U���   �E�;Er�   �M���M�U�;U�rLw�E�;E�rB�M�;M�u\�U�;U�uT�u�3��E�RPj�j������u��}��E��U��E�;E�w,r�M�;M�w"�E�RP�U�R�E�P��1��3�E�щEȉU���U���U�} u��E��M�U���U�������E���E�M��u�} t�U�U��E�    �E�    �   �E��u:�M��u{�U��t�}�   �w!r�}� w�E��uZ�}����rQw�}��vI�*��� "   �M��t�E������E������&�U��t�E�    �E�   ���E������E�����} t�E�M��U��t�E��؋M̃� �ىEȉM̋UȉU��ẺE��E������M�������E��U��M�d�    Y_^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�EP�MQ�UR�E�P�e������E���]��������������U��=4� uj �EP�MQ�URh��,�������j �EP�MQ�URj ������]����������������������������U��j �EP�MQ�UR�EP�������]������������������U��EP�MQ�UR�EP� ����]��������������������U��EP�MQ�UR�
����]��������U��EP�MQ�UR�EP������]��������������������U��=4� uj�EP�MQ�URh���������j�EP�MQ�URj � �����]����������������������������U��j�EP�MQ�UR�EP�������]������������������U��EP�MQ�UR�EP�������]��������������������U��EP�MQ�UR�EP������]��������������������U��Q�EPj �MQ�U�R�7������E���]����������������U��EP�MQ�UR������]��������U��EP�MQ��	����]������������U��EP�MQ�UR�����]��������U��EP�MQ�UR�
����]��������U��EP�MQ�UR�
����]��������U��Q�E�    ��E����E��M���M�U�;Us�E���t�ڋE���]�����������������������U����E�    �$��E��M��9 ��   j j j j j��U��Pj j ��E�}� u����   j=h�jj�M�Q�������E��}� u����rj j �U�R�E�Pj��M��Rj j ���uj�E�P�����������=j �M�Q�R�������}�}� tj�U�R��������E�    �E����E��4���3���]����������������������������������������������������������U��j �EP�MQ�UR�����]����������������������U���H�EP�M��\����} u�E�    �M������E��L  �} t	�E�   ��E�    �M��M��}� u#h8�hpjj j=h�j�5�������u̃}� u=�#���    j j=h�h\h8��������E�����M������E���  �} t	�E�   ��E�    �E�E��}� u#h��hpjj j>h�j��������u̃}� u=�#���    j j>h�h\h���P�����E�����M������E��<  �}���w	�E�   ��E�    �U�U�}� u#h�hpjj j?h�j�"�������u̃}� u=�w"���    j j?h�h\h��������E�����M�������E��   �M���(���H�y u(�UR�EP�MQ�UR�'�����EЍM������E��x�M��(���@�HQ�UR�EP�MQ�URh  �M��(���@��  Q�M��(��P�w���� �E�}� u�E�����M��[����E���U���UȍM��E����Eȋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������������U���(�} t�E�M��} t	�E�   ��E�    �U�U�}� u#h�hpjj j^h�j�0�������u̃}� u-� ���    j j^h�hh�������3��,  �} t�}|�}$~	�E�    ��E�   �M�M��}� u#hPhpjj j_h�j��������u̃}� u-� ���    j j_h�hhP�O����3��  �E�E��E�    �M�f�f�U��E����E�j�M�Q�������t�U�f�f�E��M����M����U���-u�E���E�M�f�f�U��E����E���M���+u�U�f�f�E��M����M��} u@�U�R���������t	�E
   �&�E����xt�U����Xu	�E   ��E   �}uC�M�Q��������u2�U����xt�M����Xu�E����E��M�f�f�U��E����E����3��u�E��M�Q�Y������E��}��t�V�U���A|	�E���Z~�M���a|9�U���z0�E���a|�M���z�U��� �U���E��E܋M܃�7�M���h�U�;Ur�^�E���E�M�;M�r�U�;U�u���3��u9U�w�E��EE��E���M���M�} u��U�f�f�E��M����M��*����U����U��E��u�} t�M�M��E�    �f�U��u*�E��uV�M��t	�}�   �w�U��u=�}����v4���� "   �E��t	�E�������M��t	�E�   ���E�����} t�U�E���M��t�U��ډU�E��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�:�����]����������������������U��j�EP�MQ�UR�
�����]����������������������U��j �EP�MQ�UR�������]����������������������U��j�EP�MQ�UR������]����������������������U��� �} u#hl�hpjj jdh�ej���������u̋M�M��U�R�:�����E��E��H��   u&�"��� 	   �U��B�� �M��A���  �r  �/�U��B��@t$����� "   �M��Q�� �E��P���  �A  �M��Q��tJ�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J���  ��  �E��H���U��J�E��H���U��J�E��@    �E�    �M�M��U��B%  uC����    �� �9E�t����    ���9E�u�E�P�������u�M�Q�N�����U��B%  �  �M��U��+By&h`fhpjj h�   h�ej�T�������u̋U��E��
+H�M�U��B���M���U��B���M��A�}� ~�U�R�E��HQ�U�R�������E��s�}��t!�}��t�E����M������P��M���E���U��B�� t9jj j �M�Q�������E��U�U�#U���u�E��H�� �U��J���  �c�E%��  �M��Qf��*�E�   �E%��  f�E�M�Q�U�R�E�P��������E��M�;M�t�U��B�� �M��A���  ��E%��  ��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U������3ŉE��N@  f�E�M�    �U�B    �E�@    ��M���M�U���U�} vt�E��M��P�U�@�E��MQ�o������UR�c������E�P�MQ�7������UR�G������E��M��E�    �E�    �U�R�EP�������t����M�y uB�U�B���M�A�U�B���M���M�A�U����M��U��f�U�뵋E�H�� �  u�UR������f�E�f��f�E��؋Mf�U�f�Q
�M�3��������]�������������������������������������������������������������������������������������������������U��j�hd�    P��pVW���3�P�E�d�    �EP�M��K����E�    �} t�M�U��} t	�E�   ��E�    �E�E��}� u#h�hpjj jchj�,�������u̃}� uN����    j jchh|h��������E�    �E�    �E������M�������E��U��P  �} t�}|�}$~	�E�    ��E�   �U܉U؃}� u#hPhpjj jdhj��������u̃}� uN�����    j jdhh|hP�*�����E�    �E�    �E������M��R����E��U��  �M�M��E�    �E�    �U�f�f�E��M���M�j�U�R�5������t�E�f�f�M��U���U����E���-u�M���M�U�f�f�E��M���M���U���+u�E�f�f�M��U���U�} |�}t�}$~8�} t�E�M��E�    �E�    �E������M��x����E��U���  �F�} u@�U�R�V�������t	�E
   �&�E����xt�U����Xu	�E   ��E   �}uC�M�Q��������u2�U����xt�M����Xu�E���E�M�f�f�U��E���E�E�RPj�j������EĉU��M�Q�������E�}��t�Y�U���A|	�E���Z~�M���a|9�U���z0�E���a|�M���z�U��� �U���E��EԋMԃ�7�M���   �U�;Ur�   �E���E�M�;M�rLw�U�;U�rB�E�;E�u\�M�;M�uT�u�3��E�RPj�j������u��}��E��U��U�;U�w,r�E�;E�w"�E�RP�M�Q�U�R����3�E�щẺU���U���U�} u��E�f�f�M��U���U�������E���E�M��u�} t�U�U��E�    �E�    �   �E��u:�M��u{�U��t�}�   �w!r�}� w�E��uZ�}����rQw�}��vI�v��� "   �M��t�E������E������&�U��t�E�    �E�   ���E������E�����} t�E�M��U��t�E��؋MЃ� �ىẺMЋỦU��EЉE��E������M������E��U��M�d�    Y_^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    j j j j j��EPj j ��E��}� u��P����������   h�  h�j�M�Q��������E��}� u���   j j �U�R�E�Pj��MQj j ���u!��P�B�����j�U�R���������X�E�    �E�P�MQ�U�R�E�P�������} t"�}� t�M�+M��U�J�M��	�U�    j�E�P�������E���]������������������������������������������������������������������������U��=4� uj �EP�MQ�URh����������j �EP�MQ�URj �������]����������������������������U��j �EP�MQ�UR�EP������]������������������U��EP�MQ�UR�EP�u�����]��������������������U��EP�MQ�UR������]��������U��EP�MQ�UR�EP�%�����]��������������������U��=4� uj�EP�MQ�URh����������j�EP�MQ�URj �������]����������������������������U��j�EP�MQ�UR�EP������]������������������U��EP�MQ�UR�EP�a�����]��������������������U��EP�MQ�UR�EP�1�����]��������������������U��j �EP�MQ������]����������U��EP�MQ�UR�-�����]��������U��EP�MQ�������]������������U��EP�MQ�UR�������]��������U��EP�MQ�UR������]��������U��EP�MQ�UR�������]��������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_���������������������������������U���\���3ŉE��E�E��MQ�M��,����} t�U�E��} t	�E�   ��E�    �MȉMă}� u#h�hpjj jDh�j��������u̃}� u;�i
���    j jDh�h,h���������]��M�������E��B  �M�������t/�M������ �xt~�M�����Pj�M��R�������E��j�E��Q�M����P�O������Eԃ}� t�U����U�뗍M����P�E�P�M�Q�������E܃} t�U܋E�B�M��U܋�E؋M؁�@  t���]̃} t�U�E��p�M؁�   t.�U����-u������]��	����]��A	��� "   �7�M؁�   t#�U��B��������Dz���]��	��� "   �	�E��@�]��E��]��M������E��M�3��K�����]�������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�U�����]����������U���0V�E�    �E�    �} t	�E�   ��E�    �E܉E؃}� u#hDhpjj jShpj��������u̃}� u.�����    j jShph�hD�" ��������  �U��E�}� tj=�M�Q��������E��}� t�U�;U�u�y���    ����A  �E�+E�=�  |#h�hpjj jehpj���������u�h�  �U���R������=�  r#h0hpjj jfhpj��������u̋M��Q��u	�E�   ��E�    �EԉE� �;�u� �R��  ��� ��= � ��   �} t*�=$� t!�	����t����    ����X  �   �}� t3��F  �   �= � u7h�   h�jj�������� ��= � u����  � ��     �=$� u8h�   h�jj贻�����$��=$� u�����  �$��    � ��U��}� u23�u&h�hpjj h�   hpj�Q�������u̃���  �U�+U�R�E�P�0  ���E��}� ��   �M��9 ��   j�U��E���Q�������}� ti�	�U����U��E��M��<� t�U��E��M��u��L����ց}����?s2h�   h�jj�U�R� �P�y�����E��}� t	�M�� ���U��E��M���U�    �   �}� ��   �}� }�E��؉E��M���;M�|;�U��������?s-h�   h�j�E���Pj� �Q�������E��}� u����P  �U��E��M���U��E��D�    �M�    �U�� ��j�E�P�~������M�    3��  �} ��   h  h�jj�U�R���������P�������E�}� ��   j h  hph�h �E�P�M�Q��������P�U�R������P�(������E�+E�E�E�M�� �U���U�}� t	�E�    ��E�EЋM�Q�U�R�\��u�E������}��u�^��� *   j�E�P�������}� tj�M�Q�v������U�    �E�^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    �E�E��} u3���   �M���U�E����E��}� t�M���M���h�  h�jj�U��R�������E��E��E�}� u
j	��������M�M��U��: ��   �E��Q���������E�h�  h�jj�U�R�9������M���U��: t7j h�  hph�h��E��Q�U�R�E��Q�����P�S������U����U��E����E��k����M��    �E��]������������������������������������������������������������������������������U��Q� ��E��	�M����M��U��: tK�EP�M��R�EP�s�������u/�M���E���=t�U���M���u�E�+ ����뤋E�+ ����؋�]�������������������������������������U��=4� u�EP�MQ�UR��������j �EP�MQ�UR�-����]���������������������U���H�EP�M�������} u�E�    �M������E��q  �} t	�E�   ��E�    �M��M��}� u#hhpjj j?h@j襸������u̃}� u=������    j j?h@h�h�H������E�����M��~����E���  �} t	�E�   ��E�    �E�E��}� u#h�hpjj j@h@j��������u̃}� u=�r����    j j@h@h�h���������E�����M�������E��a  �}���w	�E�   ��E�    �U�U�}� u#hLhpjj jAh@j蒷������u̃}� u=������    j jAh@h�hL�5������E�����M��k����E���   �M��d����   �� ���    u0�M��H��P�EP�MQ�UR�r������EЍM������E��   �M����� �HQ�UR�EP�MQ�URh  �M������ �   �� ���   R�M�����P������� �E�}� u�����    �E�����M������E���E���EȍM������Eȋ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���E��0}����
  �M��:}�E��0��  �U���  ��  �E=`  }�����  �M��j  }�E-`  �  �U���  }����  �E=�  }�E-�  �  �M��f	  }����w  �U��p	  }�E-f	  �]  �E=�	  }����J  �M���	  }�E-�	  �0  �U��f
  }����  �E=p
  }�E-f
  �  �M���
  }�����  �U���
  }�E-�
  ��  �E=f  }�����  �M��p  }�E-f  �  �U��f  }����  �E=p  }�E-f  �{  �M���  }����g  �U���  }�E-�  �M  �E=f  }����:  �M��p  }�E-f  �   �U��P  }����  �E=Z  }�E-P  ��   �M���  }�����   �U���  }�E-�  ��   �E=   }����   �M��*  }�E-   �   �U��@  }����   �E=J  }�E-@  �n�M���  }����]�U���  }�E-�  �F�E=  }����6�M��  }�E-  ������U���  }�E-�  ����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���X���3ŉE��E�E��MQ�M��|����} t�U�E��} t	�E�   ��E�    �MЉMԃ}� u#h�hpjj jGh�j�d�������u̃}� u;�����    j jGh�hTh����������]��M��?����E���   j�E��Q�J�������t�U����U����M�����P�E�P�M�Q�x������E܃} t�U܋B�M��A�E��M܋�U؋E�%@  t���]ȃ} t�M�U��n�E�%�   t.�M����-u������]��	����]������� "   �6�E�%   t#�M��A��������Dz���]������ "   �	�U��B�]��E��]��M��A����E��M�3��������]��������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�H�����]����������U���(���3ŉE��E�    �EPj j j j �MQ�U�R�E�P������ �E�M��t�U��   �U��E�    �E�    �F�E�P�M�Q��������E�U��u�}�u�E��   �E�M��u�}�u�U��   �U�E�M��U�+U�E�P�M�U܉Q�E��A�E�M�3��y�����]���������������������������������������������������������U��j �EP�MQ�������]����������U���4�EP�M������} t	�E�   ��E�    �M��M�}� u#hlhpjj j:h�j��������u̃}� u=�W����    j j:h�h�hl�������E�    �M�������E���   �M�������@�x u#�MQ�UR�6������E�M������E���   �	�E���E�Mf�f�U��E���t|�M������H�U��D��tS�M���M�U���u�E�    �M��F����E��j�M����U��9Mu�M���M�M������E��@��U�9Uu��h����E�9Eu�M�M��M�������E���E�    �M�������E܋�]�������������������������������������������������������������������������������������������������������U���(���3ŉE��E�    �EPj j j j �MQ�U�R�E�P������ �E�M��t�U��   �U��E�    �E�    �F�E�P�M�Q�������E�U��u�}�u�E��   �E�M��u�}�u�U��   �U�E�M��U�+U���E�P�M�U܉Q�E��A�E�M�3��G�����]������������������������������������������������������̃=@�r_�D$�����fn��p� ۋT$�   ���#���+��o
f��ft�ft�f��f��#�u����������f~�3�:E��3��D$S�����T$��   t�
��:�tY��tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u!% �t�% u��   �u�^_[3�ÍB�[ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��������������������������������������������������������������������������������������U������3ŉE��EPj j j �MQ�UR�EP�M�Q������ �E�UR�E�P�������E�}�u	�M���M�E�M�3��)�����]�����������������������������������������U���   ���3ŉE��E��E�3�f�M�ǅl���   �E�    �E�    �E�    ǅp���    �E�    ǅ|���    �E�    �E�    �E�    �E�    3�f�U�3�f�E��E�    �E�    �}$ tǅh���   �
ǅh���    ��h�����\�����\��� u#h�hpjj j~hj�V�������u̃�\��� u-�����    j j~hhh��������3���  �E�E̋M̉M��	�Ũ��ŰE���� t!�U����	t�M����
t�E����u�Ƀ}�
�N  �U�f�f�EЋM̃��M̋Uȉ�`�����`����   ��`����$�\��MЃ�1|�UЃ�9�E�   �Ẽ��E��   �MЋU$����   ��;�u	�E�   �a�EЉ�t�����t���+t��t���-t#��t���0t�*�E�   �1�E�   3�f�M��"�E�   � �  f�U���E�
   �Ẽ��E��e  �E�   �MЃ�1|�UЃ�9�E�   �Ẽ��E��|�MЋU$����   ��;�u	�E�   �[�EЉE��M���+�M��}�:w5�U������$����E�   �+�E�   �"�M̃��M��E�   ��E�
   �Ũ��U��  �EЃ�1|�MЃ�9�E�   �Ũ��U��L�EЋM$����   ��
;�u	�E�   �+�UЉ�T�����T���0t�	�E�   ��E�
   �E��E��D  �E�   ��M�f�f�UЋẼ��E��MЃ�0|:�UЃ�91�}�s �E����E��MЃ�0�U��
�E����E��	�M����M���UЋE$����   ��;�u	�E�   �R�MЉM��U���+�U��}�:w,�E�����$�؆�E�   �"�Ũ��U��E�   ��E�
   �Ẽ��E��m  �E�   �E�   �}� u)��M�f�f�UЋẼ��E��MЃ�0u�U����U�����E�f�f�MЋŨ��U��EЃ�0|8�MЃ�9/�}�s'�U����U��EЃ�0�M���U����U��E����E���MЉM��U���+�U��}�:w,�E���,��$� ��E�   �"�Ũ��U��E�   ��E�
   �Ẽ��E��  �E�   �MЃ�0|�UЃ�9�E�   �Ẽ��E���E�
   �M��M��F  �Ũ��U��EЃ�1|�MЃ�9�E�	   �Ũ��U��Y�EЉ�x�����x���+t0��x���-t��x���0t�%�E�   �)�E�   ǅl���������E�   ��E�
   �M��M��  ǅp���   ��U�f�f�EЋM̃��M��UЃ�0u���EЃ�1|�MЃ�9�E�	   �Ũ��U���E�
   �Ẽ��E��X  �MЃ�1|�UЃ�9�E�	   �Ẽ��E��+�MЉ�X�����X���0t�	�E�   ��E�
   �U��U��  ǅp���   �E�    ��E�f�f�MЋŨ��U��EЃ�0|,�MЃ�9#kU�
�EЍLЉM��}�P  ~	�E�Q  �븋U��U���E�f�f�MЋŨ��U��EЃ�0|�MЃ�9���E�
   �Ũ��U��h�}  tR�Ẽ��E��MЉ�d�����d���+t��d���-t��E�   ǅl���������E�   ��E�
   �U��U���E�
   �Ẽ��E������M�Ủ�}� �`  �}� �V  ��|��� �I  �}�vF�   k��T���|�   k��T����   k��T��E�   �U����U��E����E��}� ��   �M����M��	�U����U��E����u�U����U��E����E��ٍM�Q�U�R�E�P��������l��� }�M��ىM��U�U��U���p��� u	�E�E�E��}� u	�M�+M�M��}�P  ~	�E�   �E�}�����}ǅ|���   �0�UR�E�P�M�Q������f�U�f�U��E։E��MډM�f�U�f�U��3�f�E�3�f�M��UĉU��E��E��}� u$3�f�M�3�f�U��EĉE��M��M��U����U��Y�}� t(��  f�E��E�   ��E�    3�f�M��U����U��+��|��� t"3�f�E�3�f�M��UĉU��E��E��M����M��Uf�E�f��M�U��Q�E�M��H�U��E�ЋMf�Q
�E��M�3�������]ÍI ~�~h�����ہɂf��!���A/8S  �������  �w�n���  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������% �%�%�%�%�%�%�%�% �%$�%(�%,�%0�%4�%8�%<�%@�%D�%H�%L�%P�%T�%X�%\�%`�%d�%h�%l�%p�%t�%x�%|�%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��%��% �%�%�%�%�%�%�%�% �%$�%(�%,�%0�%4�%8�%<�%@�%D�%H�%L�%P�%T�%X�%\���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋T$�B�� ���3��y�����N�z��������������������̋T$�B�� ���3��I����0O�J��������������������̋T$�B������3������N���������������������̋T$�B������3������J�3��߀���`L���������������������������̋T$�B������3�詀���J�3�蟀����L頢�������������������������̋T$�B�� ���3��i�����M�j��������������������̋T$�B������3��9����pN�:��������������������̋T$�B������3��	����J�3������PM� ��������������������������̋M��s���M���鄝���T$�B�J�3������S麡�������������������̋M��es���T$�B�J�3�����lS酡���������������j8h���E�P�E�P�o����ËT$�B�J�3��D����R�E���������������̍M�����h���E�P�mj����ËT$�B�J�3������S������������������������������̍M�飗���T$�B�J�3���~���<S�Š���������������h�   h���E�P�E�P�h����ËT$�B�J�3��~���S邠����������������������������h�   h���E�P�E�P�kh����ËT$�B�J�3��1~����R�2����������������������������̍M��>m���T$�B�J�3���}���J�3���}����Z����������������������̍M�铖���T$�B�J�3��}����W鵟��������������̍M��c����T$�B�J�3��}���tY酟��������������̍M��3����T$�B�J�3��T}���xZ�U���������������̋M��q���T$�B�J�3��$}���TU�%���������������̋M���p���T$�B�J�3���|���pX�����������������̋M��p���T$�B�J�3���|����Y�Ş��������������̍�`����GZ���M���k����p����4Z���M���k���T$�B��0���3��s|���J�3��i|����X�j�������������������������������������h  h`��E�P�E�P�Kf����ËE����   �e���M��զ��ËT$�B�J�3���{��� U��������������������������������������hD  h`��E�P�E�P��e����ËE����   �e���M��e���ËT$�B�J�3��{���<X鉝�����������������������������������h�   h`��E�P�E�P�ke����ËE����   �e���M������ËT$�B�J�3��{����Y������������������������������������̍�\����X���M��j����`����tX���M�� j���T$�B��`���3��z���J�3��z���|W骜�����������������������������������̍�P����X���M��i����T����X���M��i���T$�B��T���3��Cz���J�3��9z����W�:������������������������������������̍M��>i���M��6i���T$�B��X���3���y���J�3���y���0W����������������������������̋T$�B��l���3��y���J�3��y���DZ頛�������������������������̍M��W���M��h���M��
W���M��h���T$�B��L���3��Iy���J�3��?y���@Y�@��������������������������̍M������T$�B�J�3��y���T����������������̍M�鰣���M�髑���T$�B�J�3���x���LT�͚�����������������������jJh���E�P�E�P�b�����jKh���E�P�E�P�b�����jLh���E�P�E�P�b�����jMh���E�P�E�P�vb�����jOh���E�P�E�P�^b����ËT$�B�J�3��$x���xT�%�����������������������������������������������̍M��U���T$�B�J�3���w���J�3���w����U�˙��������������������̍M��JU���T$�B�J�3��w���J�3��w���V鋙��������������������̍M��
U���T$�B�J�3��Tw���J�3��Jw���8V�K���������������������̍M���T���T$�B�J�3��w���J�3��
w���hV����������������������̍M��T���T$�B�J�3���v���J�3���v����V�˘��������������������̍M��JT���T$�B�J�3��v���J�3��v����V鋘��������������������̍M��
T���T$�B�J�3��Tv���J�3��Jv����V�K���������������������̍�H�����S���M��Se����|����He���M��@e����`����S���T$�B��@���3���u���J�3���u���|U�ߗ������������������������̍�p����WS���M���d���T$�B��d���3��u���J�3��u����X鍗����������������������̍M��
S���M��+����T$�B�J�3��Lu����T�M�����������������������̍M��^d���T$�B�J�3��u���J�3��
u���������������������������̍M��d���T$�B�J�3���t���J�3���t���Ѓ�˖��������������������̍M���c���T$�B�J�3��t���J�3��t���0�鋖��������������������̍M��c���T$�B�J�3��Tt���J�3��Jt������K���������������������̍M�&Z���M�Z���M��Z���M��Z���M��Z���M��IZ���M���Y���T$�B�J�3���s�������������������������������������̍M�!b���M�b���M��b���M��	b���M��b���M��HO���M���a���T$�B�J�3��ts�����u�������������������������������̋EP�E�P�^����ËT$�B�J�3��+s���@��,����������������������̋EP�E�P�V^����ËT$�B�J�3���r���������������������������̍M�铋���T$�B�J�3��r�����鵔��������������̍M��c����T$�B�J�3��r���xp酔��������������̍M��3����T$�B�J�3��Tr���w�U���������������̍M������T$�B�J�3��$r���4h�%���������������̍M��ӊ���T$�B�J�3���q���@^�����������������̍M�飊���T$�B�J�3���q���^�œ��������������̍M��s����T$�B�J�3��q����w镓��������������̍M��C����T$�B�J�3��dq����h�e���������������̍M������T$�B�J�3��4q����y�5���������������̍M������T$�B�J�3��q����j����������������̍M�鳉���T$�B�J�3���p����}�Ւ��������������̍M�郉���T$�B�J�3��p����l饒��������������̍M��S����T$�B�J�3��tp���p�u���������������̍M��#����T$�B�J�3��Dp����~�E���������������̍M������T$�B�J�3��p���$n����������������̍M��È���T$�B�J�3���o����m����������������̍M�铈���T$�B�J�3��o����s鵑��������������̍M��c����T$�B�J�3��o����d酑��������������̍M��3����T$�B�J�3��To���u�U���������������̍M������T$�B�J�3��$o���8f�%���������������̍M��Ӈ���T$�B�J�3���n���v�����������������̍M�飇���T$�B�J�3���n���<g�Ő��������������̍M��s����T$�B�J�3��n���d�镐��������������̍M��C����T$�B�J�3��dn���p�e���������������̍M������T$�B�J�3��4n������5���������������̍M������T$�B�J�3��n���Hp����������������̋M���R���T$�B�J�3���m���(~�Տ��������������̋M��R���T$�B�J�3��m����l饏��������������̋M��U���T$�B�J�3��tm���P{�u���������������̋M��*M���T$�B�J�3��Dm���p^�E���������������̋M��s����T$�B�J�3��m��� �����������������̋M���}���T$�B�J�3���l���������������������̋M���P���T$�B�J�3��l����{鵎��������������̋M��P���T$�B�J�3��l���@|酎��������������̋M��mP���T$�B�J�3��Tl���|�U���������������̋M��=P���T$�B�J�3��$l����{�%���������������̋M��P���T$�B�J�3���k����{�����������������̋M��U���T$�B�J�3���k����^�ō��������������̋M��\U���T$�B�J�3��k���`_镍��������������̋M��,U���T$�B�J�3��dk���0_�e���������������̋M���T���T$�B�J�3��4k��� _�5���������������̋M���T���T$�B�J�3��k����^����������������̋M��Qm���T$�B�J�3���j����\�Ռ��������������̋M��!m���T$�B�J�3��j���@\饌��������������̋M��U^���T$�B�J�3��tj���@v�u���������������̋M��%^���T$�B�J�3��Dj���lg�E���������������̋M��=R���T$�B�J�3��j����]����������������̋M��R���T$�B�J�3���i���(]����������������̋M��x���T$�B�J�3��i���8w鵋��������������̋M���w���T$�B�J�3��i���dh酋��������������̋M��5]���T$�B�J�3��Ti����w�U���������������̋M��]���T$�B�J�3��$i���i�%���������������̋M���\���T$�B�J�3���h����y�����������������̋M��\���T$�B�J�3���h����j�Ŋ��������������̋M��u\���T$�B�J�3��h����p镊��������������̋M��E\���T$�B�J�3��dh���b�e���������������̋M��\���T$�B�J�3��4h���t�5���������������̋M���[���T$�B�J�3��h���4e����������������̋M��[���T$�B�J�3���g���<u�Չ��������������̋M��[���T$�B�J�3��g���hf饉��������������̋M��<����T$�B�J�3��tg�����u���������������̋M������T$�B�J�3��Dg���Tn�E���������������̋M���Z���M���霏���T$�B�J�3��	g������
��������������������̋M��Z���M����\����T$�B�J�3���f����`�ʈ�������������������̍M��L���T$�B�J�3��f�����镈��������������̍M���L���T$�B�J�3��df������e���������������̍M��T���T$�B�J�3��4f���@��5���������������̍M���A���T$�B�J�3��f���p�����������������̍M���K���T$�B�J�3���e���`��Շ��������������̍M��!T���T$�B�J�3��e����饇��������������̋T$�B�J�3��|e���(}�}�����������������������̋T$�B�J�3��Le���H`�M�����������������������̍�`�����B���M��kU����p����B���M��@T���T$�B��0���3���d���J�3���d����t�������������������������������������̍�`����WB���M��kq����p����DB���M���S���T$�B��0���3��d���J�3��yd����e�z�������������������������������������h^  hЕ�E�P�E�P�[N����ËE����   �e���M�����ËT$�B�J�3��d����\�	������������������������������������hs  hЕ�E�P�E�P��M����ËE����   �e���M��u���ËT$�B�J�3��c����\际�����������������������������������jCh ��E�P�E�P�~M����ËEЃ��   �e���M��vR��ËEЃ��   �e����|�������ËT$�B�J�3��c���J�3��c���hv����������������������������������jCh ��E�P�E�P��L����ËEЃ��   �e���M���Q��ËEЃ��   �e����|����\���ËT$�B�J�3��b���J�3��ub����g�v���������������������������������hO  hЕ�E�P�E�P�[L����ËE����   �e���M�����ËT$�B�J�3��b����]�	������������������������������������hl
  hЕ�E�P�E�P��K����ËE����   �e���M��u���ËT$�B�J�3��a���h]陃�����������������������������������jMh���E�P�E�P�~K����ËE����   �e���M�����ËT$�B�J�3��+a���xw�,�����������������������jMh���E�P�E�P�K����ËE����   �e���M�騋��ËT$�B�J�3���`����h�̂����������������������h�  h��E�P�E�P�J����ËE����   �e���M��E���ËT$�B�J�3��h`���x�i������������������������������������h�  h��E�P�E�P�KJ����ËE����   �e���M��Պ��ËT$�B�J�3���_���Hi��������������������������������������h�  h��E�P�E�P��I����ËE����   �e���M��e���ËT$�B�J�3��_����y鉁�����������������������������������h�  h��E�P�E�P�kI����ËE����   �e���M������ËT$�B�J�3��_���$k�������������������������������������h(  h��E�P�E�P��H����ËE����   �e���M�酉��ËT$�B�J�3��^���<驀�����������������������������������h(  h��E�P�E�P�H����ËE����   �e���M�����ËT$�B�J�3��8^����~�9������������������������������������h(  h��E�P�E�P�H����ËE����   �e���M�饈��ËT$�B�J�3���]����m�������������������������������������h(  h��E�P�E�P�G����ËE����   �e���M��5���ËT$�B�J�3��X]���|m�Y�����������������������������������h  h`��E�P�E�P�;G����ËE����   �e���M��Ň��ËT$�B�J�3���\����p��~�����������������������������������h  h`��E�P�E�P��F����ËE����   �e���M��U���ËT$�B�J�3��x\����a�y~�����������������������������������hD  h`��E�P�E�P�[F����ËE����   �e���M�����ËT$�B�J�3��\����s�	~�����������������������������������hD  h`��E�P�E�P��E����ËE����   �e���M��u���ËT$�B�J�3��[��� e�}�����������������������������������h�   h`��E�P�E�P�{E����ËE����   �e���M�����ËT$�B�J�3��([���|u�)}�����������������������������������h�   h`��E�P�E�P�E����ËE����   �e���M�镅��ËT$�B�J�3��Z����f�|�����������������������������������h�   h|��E�P�E�P�D����ËE����   �e���M��%���ËT$�B�J�3��HZ�����I|�����������������������������������h�   h|��E�P�E�P�+D����ËE����   �e���M�鵄��ËT$�B�J�3���Y����n��{�����������������������������������h  h|��E�P�E�P�C����ËE����   �e���M��E���ËT$�B�J�3��hY������i{�����������������������������������h|  h|��E�P�E�P�KC����ËE����   �e���M��Ճ��ËT$�B�J�3���X���4a��z����������������������������������̍�L����g6���M���G����P����T6���M���G���T$�B��P���3��X���J�3��X���s�z�����������������������������������̍�L�����5���M��G����P�����5���M��pG���T$�B��P���3��#X���J�3��X���@d�z�����������������������������������̍�0����5���M��G����4����t5���M�� G���T$�B��4���3��W���J�3��W���`s�y�����������������������������������̍�0����5���M��F����4����5���M��F���T$�B��4���3��CW���J�3��9W����d�:y�����������������������������������̍M��4���T$�B�J�3���V���4���x��������������̍M��z4���T$�B�J�3���V����o��x��������������̍M���E���M���E���T$�B��8���3��V���J�3��V����r�x�������������������������̍M��E���M��E���T$�B��8���3��9V���J�3��/V����c�0x�������������������������̍������3���������3���M��@F���M�� E���������3���M��%F��������<����h����;����|������   ��|������\����;��Í�D����;����|������   ��|������������E��Ë�|������   ��|�����������E��Ë�|������   ��|����������}E��Ë�|������   ��|��������[E��Í�d����7D���M��/D���������7;����,�����:����|����� �   ��|���ߍ�P�����:��Í�8����:���T$�B��0���3��T���J�3��T����x�v���������������������������������������������������������������������������������������������������������������̍������1���������1���M���`���M��0C���������1���M��`��������/����h����:B����|������   ��|������\����B��Í�D����B����|������   ��|�����������A`��Ë�|������   ��|�����������`��Ë�|������   ��|�����������_��Ë�|������   ��|���������_��Í�d����GB���M��?B���������.����,����\A����|����� �   ��|���ߍ�P����;A��Í�8����/A���T$�B��0���3��R���J�3��R����i�t���������������������������������������������������������������������������������������������������������������̋T$�B�J�3��R���J�3��R����~�t������������̋T$�B�J�3���Q���J�3���Q���8m��s������������̋T$�B��l���3��Q���J�3��Q����u�s�������������������������̋T$�B��l���3��yQ���J�3��oQ���g�ps�������������������������̋T$�B�J�3��<Q���@��=s����������������������̋T$�B�J�3��Q����n�s����������������������̍M��gy���T$�B�J�3���P������r��������������̍M��7y���T$�B�J�3��P���ha�r��������������̍M��*.���M���@���M��.���M��?���T$�B��L���3��YP���J�3��OP����t�Pr�������������������������̍M���-���M���\���M��-���M��F?���T$�B��L���3���O���J�3���O���f��q��������������������������jUh��E�P�E�P��9�����jVh���P���P�E�P��9�����jWh���8���P�E�P�9�����jXh���H���P�E�P�9�����jYh���(���P�E�P�r9�����jZh���@���P�E�P�W9�����j[h���0���P�E�P�<9�����j\h���|���P�E�P�!9�����j]h���l���P�E�P�9�����j^h���\���P�E�P��8�����j_h���L���P�E�P��8�����j`h���<���P�E�P�8�����jbh���,���P�E�P�8����ËT$�B��,���3��]N���l[�^p��������������������������������������������������������������������������������������������������������j-h��E�P�E�P��7�����j.h���P���P�E�P��7�����j/h���8���P�E�P��7�����j0h���H���P�E�P�7�����j1h���(���P�E�P�7�����j2h���@���P�E�P�w7�����j3h���0���P�E�P�\7�����j4h���|���P�E�P�A7�����j5h���l���P�E�P�&7�����j6h���\���P�E�P�7�����j7h���L���P�E�P��6�����j8h���<���P�E�P��6�����j:h���,���P�E�P�6����ËT$�B��,���3��}L����Z�~n�������������������������������������������������������������������������������������������������������̍M�Q2���M�I2���T$�B�J�3���K����}��m����������������������̍M�'���M�x'���T$�B�J�3��K����`�m����������������������̍M��1���T$�B�J�3��tK����}�um��������������̍M�'���T$�B�J�3��DK���|l�Em��������������̍M$�v;���������(����t����(���M��@:���M��P;���M��H;���������0����$�����0���������0����������0����������0���������0���������0���������0���� ����0���T$�B��t���3��J���J�3��vJ����z�wl����������������������������������������������������������������̍M$��V���������'����t����'���M��@9���M���V���M��V��������X8����$����M8��������B8���������78���������,8���������!8���������8���������8���� ���� 8���T$�B��t���3��I���J�3��vI����k�wk����������������������������������������������������������������̍M��^8���T$�B�J�3��I���J�3��
I���Px�k��������������������̍M��8���T$�B�J�3���H���J�3���H����x��j��������������������̍M���7���T$�B�J�3��H���J�3��H���|i�j��������������������̍M��7���T$�B�J�3��TH���J�3��JH����i�Kj��������������������̍M���%���T$�B�J�3��H���J�3��
H���pq�j��������������������̍M��%���T$�B�J�3���G���J�3���G����q��i��������������������̍M��J%���T$�B�J�3��G���J�3��G����q�i��������������������̍M��
%���T$�B�J�3��TG���J�3��JG��� r�Ki��������������������̍M���$���T$�B�J�3��G���J�3��
G����r�i��������������������̍M��$���T$�B�J�3���F���J�3���F���0r��h��������������������̍M��J$���T$�B�J�3��F���J�3��F���`r�h��������������������̍�H����$���M��6����|����6���M��6����`�����#���T$�B��@���3��(F���J�3��F���q�h������������������������̍M��#���T$�B�J�3���E���J�3���E����b��g��������������������̍M��Z#���T$�B�J�3��E���J�3��E����b�g��������������������̍M��#���T$�B�J�3��dE���J�3��ZE����b�[g��������������������̍M���"���T$�B�J�3��$E���J�3��E���,c�g��������������������̍M��"���T$�B�J�3���D���J�3���D����c��f��������������������̍M��Z"���T$�B�J�3��D���J�3��D���\c�f��������������������̍M��"���T$�B�J�3��dD���J�3��ZD����c�[f��������������������̍�H�����!���M���P����|�����P���M���P����`����!���T$�B��@���3���C���J�3���C���@b��e������������������������̍M��j!���T$�B�J�3��C�����e��������������̍M��:!���T$�B�J�3��C����o�e��������������̍M��
!���T$�B�J�3��TC������Ue��������������̍M��� ���T$�B�J�3��$C���Xo�%e��������������̍M�� ���T$�B�J�3���B���t���d��������������̍M��z ���T$�B�J�3���B���(o��d��������������̍M��J ���T$�B�J�3��B���Ԁ�d��������������̍M�� ���T$�B�J�3��dB����o�ed��������������̍M������M��2���T$�B�J�3��,B���J�3��"B���pz�#d����������������������������̍M�����M��>2���T$�B�J�3���A���J�3���A���4z��c����������������������������̍M��J���M��^N���T$�B�J�3��A���J�3��A����k�c����������������������������̍M������M��N���T$�B�J�3��<A���J�3��2A���`k�3c����������������������������̍�p�������M��K1���T$�B��d���3���@���J�3���@���@t��b����������������������̍�p����W���M��kM���T$�B��d���3��@���J�3��@���le�b����������������������̍M��&M���M���.���T$�B�J�3��L@���J�3��B@���L��Cb����������������������������̍M���L���M��y.���T$�B�J�3���?���J�3���?����a��a����������������������������̍M��0���M��%���M��%���T$�B�J�3��?���J�3��?����v�a��������������������̍M��6L���M���-���M���-���T$�B�J�3��T?���J�3��J?��� h�Ka��������������������̋E����   �e���M��N.��ËT$�B�J�3��?���J�3���>���\��`�������������������̍M,��$���M ��$���M�%���M�	%���M��%����p����$���M���$����|�����$����d����$���M���$���T$�B��l���3��p>���h|�q`������������������������������������������̍M,�,���M �,���M�����M�����M�������p����v,���M������|��������d����X,���M�����T$�B��l���3���=����_��_������������������������������������������̍M�:���M�:���M��:���M��:���M��:���M��$���M��|:���T$�B�J�3��T=���L��U_������������������������������̍M���U���T$�B�J�3��=������_��������������̍M���U���T$�B�J�3���<���8���^��������������̍M��U���T$�B�J�3��<�����^��������������̍M��cU���T$�B�J�3��<�����^��������������̍M��3U���T$�B�J�3��T<������U^��������������̍M��U���T$�B�J�3��$<�����%^��������������̍M���T���T$�B�J�3���;���x���]��������������̍M��T���T$�B�J�3���;�������]��������������̋M�� ���T$�B�J�3��;���<��]��������������̋M��QA���T$�B�J�3��d;���p��e]��������������̋M��/���T$�B�J�3��4;���̇�5]��������������̋M��\I���T$�B�J�3��;���Ĉ�]��������������̋M��.���T$�B�J�3���:���h���\��������������̋M��.���T$�B�J�3��:���D��\��������������̋M��<`���T$�B�J�3��t:������u\��������������̋M��%.���M�����b���T$�B�J�3��9:������:\�������������������̍M��,7���T$�B�J�3��:������\��������������̍M��!���T$�B�J�3���9���$���[��������������̍M���6���T$�B�J�3��9���đ�[���������������jCh ��E�P�E�P�#����ËEЃ��   �e���M��(��ËEЃ��   �e����|����d��ËT$�B�J�3��/9���J�3��%9�����&[��������������������������������jMh���E�P�E�P�#����ËE����   �e���M��c��ËT$�B�J�3��8�����Z����������������������h�  h��E�P�E�P�"����ËE����   �e���M��5c��ËT$�B�J�3��X8������YZ�����������������������������������h�  h��E�P�E�P�;"����ËE����   �e���M���b��ËT$�B�J�3���7�������Y�����������������������������������h(  h��E�P�E�P��!����ËE����   �e���M��Ub��ËT$�B�J�3��x7���P��yY�����������������������������������h(  h��E�P�E�P�[!����ËE����   �e���M���a��ËT$�B�J�3��7���܍�	Y�����������������������������������h�   h|��E�P�E�P�� ����ËE����   �e���M��ua��ËT$�B�J�3��6�����X�����������������������������������h�  h|��E�P�E�P�{ ����ËE����   �e���M��a��ËT$�B�J�3��(6������)X����������������������������������̍M�����T$�B�J�3���5���H���W��������������̍������g���������\���M���$���M���$���������A���M���$������������x����2����|������   ��|������l����t2��Í�T����h2����|������   ��|�����������i$��Ë�|������   ��|�����������G$��Ë�|������   ��|������,����%$��Ë�|������   ��|�������$��Í�d�����#���M���#�������������<����1����|����� �   ��|���ߍ�`����1��Í�H����1���T$�B��@���3��_4���J�3��U4���4��VV���������������������������������������������������������������������������������������������������������������̋T$�B�J�3���3���J�3���3�������U������������̋T$�B�J�3��3���T��U����������������������̍M���[���T$�B�J�3��d3���(��eU���������������j'hа�E�P�E�P�^�����j(hа�E�P�E�P�F�����j)hа�E�P�E�P�.�����j*hа�E�P�E�P������j+hа�E�P�E�P�������j,hа�E�P�E�P�������j-hа�E�P�E�P�������j.hа��x���P�E�P�����ËT$�B��|���3��v2���T��wT����������������������������������������������������������������̍M�M���M�E���T$�B�J�3��2���(��T����������������������̍M����T$�B�J�3���1���܌��S��������������̍M$�� ���������O����t����D���M��� ���M��� ���M��� ��������.����$����.��������}.���������r.���������g.���������\.���������Q.���������F.���� ����;.���T$�B��t���3��1���J�3��1���(��S����������������������������������������������������������������̍M������T$�B�J�3��0���J�3��0���܉�R��������������������̍M�����T$�B�J�3��d0���J�3��Z0�����[R��������������������̍M������T$�B�J�3��$0�����%R��������������̍M�����T$�B�J�3���/�������Q��������������̍M��z���T$�B�J�3���/�������Q��������������̍M��J���T$�B�J�3��/�����Q��������������̍M�����M�����T$�B�J�3��\/���J�3��R/������SQ����������������������������̍M������M��V���T$�B�J�3��/���J�3��/������Q����������������������������̍M�����M���+���T$�B�J�3��.���J�3��.���`��P����������������������������̍M�����M��+���M��+���T$�B�J�3��d.���J�3��Z.���`��[P��������������������̍M,�L+���M �D+���M�M���M�E���M��=����p����!+���M��*����|��������d����+���M�����T$�B��l���3���-�������O������������������������������������������̋T$�B�J�3��-���L��O����������������������̍M��(���T$�B�J�3��T-���h��UO��������������̍M��(���T$�B�J�3��$-�����%O��������������̡������ËT$�B�J�3���,���X���N������������������������̍M��(���T$�B�J�3��,�����N��������������̍M���'���T$�B�J�3��,���8��N��������������̍M��'���T$�B�J�3��T,���h��UN�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ���������'��_^[���   ;���4����]���������������������U����   SVW��@����0   ���������e��_^[���   ;��4����]���������������������U����   SVW��@����0   ���������eI��_^[���   ;��[4����]���������������������U����   SVW��@����0   ������������_^[���   ;��4����]���������������������U����   SVW��@����0   ����������_^[���   ;��3����]���������������������U����[��]������������������U�������]������������������U����� ��]������������������U�����0H��]������������������U�����2��]������������������U�������]������������������U������G��]������������������U�칲��3��]������������������U�칼��u���]������������������U�������]������������������U����� ��]������������������U�����0G��]������������������U�����2��]������������������U�������]������������������U������F��]������������������U��������]������������������U�����@��]������������������U�����pF��]������������������U�����r��]������������������U��������]������������������U�����F��]������������������U��g������]������������������U��d����]������������������U������ ��]������������������U�����@��]������������������U�����pE��]������������������U�����r ��]������������������U��������]������������������U�����E��]������������������U����� ��]������������������U�������]������������������U�����D��]������������������U��������]������������������U����� ��]������������������U�����PD��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                           0�����    �������� � �@�����@� ���`����� �`��� ��������������P�0����                                                                                                                                                                                                                                                                                            p�������p���P�                                                                                                                                                                                                                                                                        �����    ��@���P�����@� �����������p�    �P�����    ����    ����    P�@�     ���    ����    @�0�    � �    @�0�    p�`�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �q>(r?E                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            |&�$                                                                                                                                                                                                                                                                    ^                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                P�Z       s   � ��     P�Z          � �� lP4B�h1E]P9D@ <6        c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ x u t i l i t y                               I T E R A T O R   L I S T   C O R R U P T E D !             ����#�#"l    bad locale name     t#�$�_�_    $A�A8e    c:\program files (x86)\microsoft visual studio 12.0\vc\include\xlocale                  ($�j�A8e�&VGCd            c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ x l o c a l e                                 �$�.�A8e    �$I;�A8e�&Zu@0�C3�^Qt�Y            L%7\�_�_�_�P�&        �%�'"l    :   &(M"l    h&^gG�7�_�P�&        generic     unknown error   �&�O�3�n�_�P�&        iostream    iostream stream error       $'�2?O�`wX�P�&        system  �'
M"l     �9    ios_base::badbit set        ios_base::failbit set       ios_base::eofbit set            c:\program files (x86)\microsoft visual studio 12.0\vc\include\xiosbase                 � �Q    �!�#               (!]^%-�7']W�A�>Fk�/@gVByG.[�j9            P"�6�lg=Q�>�A�[�!�/@g�o0rX�X�g            �"HF        p       ERROR: COULD NOT READ FILE      T(�,�)�h1E]P9D@ <6        Load .stl File      STL solid   Ascii stl Files Not Supported!              c:\program files\maxon\cinema 4d r13\plugins\stl_importer\source\stl_importer.cpp                   STL Importer    stl_icon.png        c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ x s t r i n g                                     c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ i s t r e a m                                 i >= 0 && i < count         c:\program files\maxon\cinema 4d r13\resource\_api\ge_dynamicarray.h                %s(%d): %s      �'�%�A8eg6VGCd�%G.|NXJ        c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ v e c t o r                               v e c t o r   i t e r a t o r   n o t   d e r e f e r e n c a b l e                 Standard C++ Libraries Out of Range         " S t a n d a r d   C + +   L i b r a r i e s   O u t   o f   R a n g e "   & &   0                     % s     s t d : : _ V e c t o r _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ V e c t o r _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < s t r u c t   t r i a n g l e >   >   > : : o p e r a t o r   *                                               " o u t   o f   r a n g e "             v e c t o r   i t e r a t o r   n o t   i n c r e m e n t a b l e                       s t d : : _ V e c t o r _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ V e c t o r _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < s t r u c t   t r i a n g l e >   >   > : : o p e r a t o r   + +                                                 string too long     invalid string position         c:\program files (x86)\microsoft visual studio 12.0\vc\include\streambuf                vector<T> too long      v e c t o r   i t e r a t o r s   i n c o m p a t i b l e               Standard C++ Libraries Invalid Argument         " S t a n d a r d   C + +   L i b r a r i e s   I n v a l i d   A r g u m e n t "   & &   0                     s t d : : _ V e c t o r _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ V e c t o r _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < s t r u c t   t r i a n g l e >   >   > : : _ C o m p a t                                             " i n v a l i d   a r g u m e n t "             s t r i n g   i t e r a t o r   n o t   d e r e f e r e n c a b l e                     s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < c h a r >   >   > : : o p e r a t o r   *                                             i n v a l i d   n u l l   p o i n t e r             bad cast    i n v a l i d   i t e r a t o r   r a n g e             FALSE   c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ x m e m o r y                                     c:\program files\maxon\cinema 4d r13\resource\_api\c4d_resource.cpp                 #   M_EDITOR        c:\program files\maxon\cinema 4d r13\resource\_api\c4d_memory.cpp               c:\program files\maxon\cinema 4d r13\resource\_api\c4d_string.cpp               no baselist      GB  MB  KB  B        �@    �(fi    c:\program files\maxon\cinema 4d r13\resource\_api\c4d_file.cpp             res                       �?        c:\program files\maxon\cinema 4d r13\resource\_api\c4d_general.h                   %s  �(�M)t    $)�_    |)Rn    c:\program files\maxon\cinema 4d r13\resource\_api\c4d_baseobject.cpp               nncnt<ncnt      nncnt==ncnt         ����MbP?        c:\program files\maxon\cinema 4d r13\resource\_api\c4d_pmain.cpp                c:\program files\maxon\cinema 4d r13\resource\_api\c4d_basebitmap.cpp               c:\program files\maxon\cinema 4d r13\resource\_api\ge_sort.cpp              c:\program files\maxon\cinema 4d r13\resource\_api\c4d_libs\lib_ngon.cpp                      �?        ������        �������    �)Xm    0*�i    �*�U    c:\program files\maxon\cinema 4d r13\resource\_api\c4d_gv\ge_mtools.cpp                 �*�i                                                                                                         	           	         	       �x     �x     �x   H   �x       �x      �x      �x     �x      �x   �  �x      �x   H   �x   H   �x      �x   ��  �x   �                                                           	   alnum   alpha   blank   cntrl   d   digit   graph   lower   print   punct   space  s   upper   w   xdigit  ?          @      z     z     ,z   H   <z       Lz      Pz      `z     pz      �z   �  �z      �z   H   �z   H   �z      �z   ��  �z   �                                                             	   �   &   ����a l n u m       a l p h a       ����b l a n k       c n t r l       d   d i g i t       g r a p h       l o w e r       p r i n t       p u n c t       s p a c e       s   u p p e r       w   x d i g i t     5            4  �������5            4  �������                   @   �                           0   @   �  �      0                                 @   �                                                        ?                                                                            <+�q"l    bad allocation      �+�k"l    �+("l    T,�Z"l    �,{O"l    -�D"l    t-8�c    bad function call       �-�s"l        regex_error(error_collate): The expression contained an invalid collating element name.                         regex_error(error_ctype): The expression contained an invalid character class name.                     regex_error(error_escape): The expression contained an invalid escaped character, or a trailing escape.                         regex_error(error_backref): The expression contained an invalid back reference.                 regex_error(error_brack): The expression contained mismatched [ and ].                  regex_error(error_paren): The expression contained mismatched ( and ).                  regex_error(error_brace): The expression contained mismatched { and }.                  regex_error(error_badbrace): The expression contained an invalid range in a { expression }.                     regex_error(error_range): The expression contained an invalid character range, such as [b-a] in most encodings.                         regex_error(error_space): There was insufficient memory to convert the expression into a finite state machine.                          regex_error(error_badrepeat): One of *?+{ was not preceded by a valid regular expression.                       regex_error(error_complexity): The complexity of an attempted match against a regular expression exceeded a pre-set level.                              regex_error(error_stack): There was insufficient memory to determine whether the regular expression could match the specified character sequence.                               regex_error(error_parse)        regex_error(error_syntax)       regex_error     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x s t r i n g                   f:\dd\vctools\crt\crtw32\stdcpp\_tolower.c          f:\dd\vctools\crt\crtw32\stdcpp\locale0.cpp         0.�u�A8e    *   C   f:\dd\vctools\crt\crtw32\stdhpp\xutility                      ��    �   0�o   D��   \��   \�R   ��  x��  x��  x�   �7   0�d	  \��   ��  ��p   ��P    �   Ȋ'   ��   �   0�   �   ��{   ��!   ��   ��   ���  �   �   4�   \�n   x�a	  \��  t�   �   Ȋ   x��  4�   x�    �   ��   x�   �'  ��@'  ��A'  Ћ?'  �5'  �'  8�E'  P�M'  h�F'  ��7'  ��'  ��Q'  Ȍ4'  ܌'  ��&'  �H'  �('  4�8'  L�O'  \�B'  t�D'  ��C'  ��G'  ��:'  ��I'  ؍6'  �='  ��;'  �9'  0�L'  H�3'  T�        f   p�d   ��e   ��q   Ď   ܎!   ��   �	   $�h   <�    L�j   \�g   t�k   ��l   ��   \�m   ȏ   \�)   ��   �    �   �&   D�(   �n   �o   0�*   H�   d�   ��   ��   ��   x�   ��s   ��t   Đu   Ԑv   �w   ��
   �y   $�'   �x   0�z   L�{   \�   ��|   t�   ��   0�   Ȋ   ��   ���   ԑ}   �~   ��   ��   �i   t�p   �   0��   L��   h��   ��   ��   ���   ��   Ē$   ��   4�"   �   ��   8��   L��   `�   l�   ��   ��r   ���   ȓ�   ܓ                                                                                                                                                                                                                                                                permission denied       file exists     no such device      filename too long       device or resource busy     io error    directory not empty     invalid argument    no space on device      no such file or directory       function not supported      no lock available       not enough memory       resource unavailable try again          cross device link       operation canceled      too many files open     permission_denied       address_in_use      address_not_available       address_family_not_supported        connection_already_in_progress          bad_file_descriptor     connection_aborted      connection_refused      connection_reset    destination_address_required        bad_address     host_unreachable    operation_in_progress       interrupted     invalid_argument    already_connected       too_many_files_open     message_size    filename_too_long       network_down    network_reset   network_unreachable     no_buffer_space     no_protocol_option      not_connected   not_a_socket    operation_not_supported     protocol_not_supported      wrong_protocol_type     timed_out   operation_would_block       address family not supported        address in use      address not available       already connected       argument list too long      argument out of domain      bad address     bad file descriptor     bad message     broken pipe     connection aborted      connection already in progress          connection refused      connection reset    destination address required        executable format error     file too large      host unreachable    identifier removed      illegal byte sequence       inappropriate io control operation          invalid seek    is a directory      message size    network down    network reset   network unreachable     no buffer space     no child process    no link     no message available        no message      no protocol option      no stream resources     no such device or address       no such process     not a directory     not a socket    not a stream    not connected   not supported   operation in progress       operation not permitted     operation not supported     operation would block       owner dead      protocol error      protocol not supported      read only file system       resource deadlock would occur       result out of range     state not recoverable       stream timeout      text file busy      timed out   too many files open in system       too many links      too many symbolic link levels       value too large     wrong protocol type         ��������                    `��x�xd�h�l�l�p�t�x�|�������                r   a   rb  wb  ab  r+  w+  a+  r+b w+b a+b Ԕ�z�zؔܔ����������$�                r   a   r b     w b     a b     r +     w +     a +     r + b       w + b       a + b                
   !   "   2   *            #   3   +                            
   !   "   2   *            #   3   +                   false   true    f:\dd\vctools\crt\crtw32\stdhpp\xlocale         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x l o c a l e                   f:\dd\vctools\crt\crtw32\stdhpp\xlocnum         f:\dd\vctools\crt\crtw32\stdcpp\locale.cpp          �.�@�A8e�&�)))�.�.)e)j))~.            �.4n�A8e�C)))�a�a�(�(_a            P/)j�A8evOo�kT]�^            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x l o c n u m                   ld  lu  Ld  Lu  %p  0123456789ABCDEFabcdef-+Xx      0123456789-+Ee      eE  pP  .   s t r i n g   s u b s c r i p t   o u t   o f   r a n g e               0123456789ABCDEFabcdef-+XxPp        f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ s t r e a m b u f                       i s t r e a m b u f _ i t e r a t o r   i s   n o t   d e r e f e r e n c a b l e                       i s t r e a m b u f _ i t e r a t o r   i s   n o t   i n c r e m e n t a b l e                         z�����8            _�B        �M�raB3G        f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x u t i l i t y                         :Sun:Sunday:Mon:Monday:Tue:Tuesday:Wed:Wednesday:Thu:Thursday:Fri:Friday:Sat:Saturday                   :Jan:January:Feb:February:Mar:March:Apr:April:May:May:Jun:June:Jul:July:Aug:August:Sep:September:Oct:October:Nov:November:Dec:December                                  : S u n : S u n d a y : M o n : M o n d a y : T u e : T u e s d a y : W e d : W e d n e s d a y : T h u : T h u r s d a y : F r i : F r i d a y : S a t : S a t u r d a y                                       : J a n : J a n u a r y : F e b : F e b r u a r y : M a r : M a r c h : A p r : A p r i l : M a y : M a y : J u n : J u n e : J u l : J u l y : A u g : A u g u s t : S e p : S e p t e m b e r : O c t : O c t o b e r : N o v : N o v e m b e r : D e c : D e c e m b e r                                                         �/uZ�A8e�(D6E+�]�H�6�N        0�!�A8e"S�Q�(�l�]k(7C        x0}%�A8e]YI,33�u�L9Z_�dXr/�a�Q            �0�]�A8e�d�$a_�:#k~L�%!'�$�a/(ED            ����`2�H�A8e    �2�+�A8e     3�i�A8e    �6>�A8e�Y    f:\dd\vctools\crt\crtw32\stdcpp\wlocale.cpp         @1U>�A8e�gQjj�i�%=$Uk�jZk�j&            �3$8�A8e�+\
\5	5Z/Z5             2?�A8eR<�i9d�E�T        �3�+�A8e/s�n(f        @4Pk�A8e�f5@�         �4�R�A8e�5�X    5�Q�A8e	b�]    L7�E�A8eNJ�<^q�2K%�0M�H�;            d5ks�A8eNJ�<^q�2K%�0M�H�;            6d9�A8eNJ�<^q�2K%�0M�H�;            �6�n�A8e�E�9:6cb)B�]N6        �1BL�A8e�%:'?''`[[7%<%#%n%[[            d7Yq�A8e5'�2�2qrgr33r            �7X6�A8e�'�>�[T+�*        $8l�A8e�:�At        �8L=�A8e�8�Dk-        �8u-�A8e�5�;    ����H9C2�A8egE�0    �;k#�A8eytsHmg�5�d�4S6�(�"            �9XY�A8eytsHmg�5�d�4S6�(�"            `:�G�A8eytsHmg�5�d�4S6�(�"            �:K�A8e5,�_Bo6i4ZC�>        0;�;�A8e�R    f:\dd\vctools\crt\crtw32\stdhpp\xloctime            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x l o c t i m e                     ! % x       f:\dd\vctools\crt\crtw32\stdhpp\locale          f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ l o c a l e                     f:\dd\vctools\crt\crtw32\stdhpp\xlocmes         f:\dd\vctools\crt\crtw32\stdhpp\xlocmon         %.0Lf   0123456789-     %b %d %H : %M : %S %Y       %m / %d / %y        :AM:am:PM:pm    %I : %M : %S %p     %H : %M     %H : %M : S     %d / %m / %y    0123456789-     0123456789ABCDEFabcdef-+Xx      0123456789-+Ee          f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x l o c m o n                   0123456789-     0123456789ABCDEFabcdef-+Xx      0123456789-+Ee      0123456789-     0123456789ABCDEFabcdef-+XxPp        $+xv    : A M : a m : P M : p m         0123456789ABCDEFabcdef-+XxPp            s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < w c h a r _ t >   >   > : : o p e r a t o r   *                                               s t r i n g   i t e r a t o r   n o t   i n c r e m e n t a b l e                       s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < w c h a r _ t >   >   > : : o p e r a t o r   + +                                             s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < u n s i g n e d   s h o r t >   >   > : : o p e r a t o r   *                                                 s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < u n s i g n e d   s h o r t >   >   > : : o p e r a t o r   + +                                                   -   +v$x+v$xv$+xv+$xv$+x+$vx+$vx$v+x+$vx$+vx+v $+v $v $+v +$v $++$ v+$ v$ v++$ v$+ v+xv$+ v$v$ +v+ $v$ ++x$v+ $v$v ++ $v$ +v                                s t r i n g   i t e r a t o r   +   o f f s e t   o u t   o f   r a n g e                       s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < w c h a r _ t >   >   > : : o p e r a t o r   + =                                             s t r i n g   i t e r a t o r s   i n c o m p a t i b l e               s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < w c h a r _ t >   >   > : : _ C o m p a t                                             s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < u n s i g n e d   s h o r t >   >   > : : o p e r a t o r   + =                                               s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < u n s i g n e d   s h o r t >   >   > : : _ C o m p a t                                               -   �;�M�A8e2%sj        f:\dd\vctools\crt\crtw32\stdcpp\xlocale.cpp         <uP�A8e�O�bdC        l<@D�A8e�n�H    �<�A�A8eA�%    ?sC�A8eW�n�S�P�f�d7>�5�N            ,=�c�A8eW�n�S�P�f�d7>�5�N            �=�F�A8eW�n�S�P�f�d7>�5�N            P>m:�A8e�e�$~o�,Is/P         �>Y5�A8e=)    0123456789-     !%x     0123456789-         s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < c h a r >   >   > : : o p e r a t o r   + +                                           s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < c h a r >   >   > : : o p e r a t o r   + =                                           s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < c h a r >   >   > : : _ C o m p a t                                                 �M(knN          �A            e��A    0123456789abcdefghijklmnopqrstuvwxyz      !

					               0123456789abcdefghijklmnopqrstuvwxyz      A)!                   p l o c - > _ M b c u r m a x   = =   1   | |   p l o c - > _ M b c u r m a x   = =   2                         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d c p p \ x m b t o w c . c                   f:\dd\vctools\crt\crtw32\stdcpp\xwcsxfrm.c          0123456789abcdefABCDEF   	

            �?  �? @F   �  �� ��= �9 �3       A      �?              �              �           ����?   ���9>   033�<              $@           ����?   ���9>   033�<           ?  � ������?�                      ?  � ������?�                         f:\dd\vctools\crt\crtw32\misc\onexit.c          ���    d s t   ! =   N U L L       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ m e m c p y _ s . c                     m e m c p y _ s         s r c   ! =   N U L L       s i z e I n B y t e s   > =   c o u n t             ,?Z/"l    Unknown exception       D?�,"l    �?H"l    �?q"l    ( s t r e a m   ! =   N U L L )         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f c l o s e . c                   f c l o s e     ( s t r   ! =   N U L L )           _ f c l o s e _ n o l o c k         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f g e t c . c                     f g e t c       (   ( _ S t r e a m - > _ f l a g   &   _ I O S T R G )   | |   (   f n   =   _ f i l e n o ( _ S t r e a m ) ,   (   ( _ t e x t m o d e _ s a f e ( f n )   = =   _ _ I O I N F O _ T M _ A N S I )   & &   ! _ t m _ u n i c o d e _ s a f e ( f n ) ) ) )                                                       g e t c     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f g e t p o s . c                     f g e t p o s       ( p o s   ! =   N U L L )               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f p u t c . c                     f p u t c       p u t c         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f s e t p o s . c                     f s e t p o s       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f s e e k i 6 4 . c                   _ f s e e k i 6 4           ( ( w h e n c e   = =   S E E K _ S E T )   | |   ( w h e n c e   = =   S E E K _ C U R )   | |   ( w h e n c e   = =   S E E K _ E N D ) )                                 s t r   ! =   N U L L       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f w r i t e . c                   f w r i t e     _ f w r i t e _ n o l o c k         ( b u f f e r   ! =   N U L L )         n u m   < =   ( S I Z E _ M A X   /   s i z e )             ( " I n c o n s i s t e n t   S t r e a m   C o u n t .   F l u s h   b e t w e e n   c o n s e c u t i v e   r e a d   a n d   w r i t e " ,   s t r e a m - > _ c n t   > =   0 )                                             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ s e t v b u f . c                     s e t v b u f       ( t y p e   = =   _ I O N B F )   | |   ( t y p e   = =   _ I O F B F )   | |   ( t y p e   = =   _ I O L B F )                         ( ( 2   < =   s i z e )   & &   ( s i z e   < =   I N T _ M A X ) )                 f:\dd\vctools\crt\crtw32\stdio\setvbuf.c            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ u n g e t c . c                   u n g e t c     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ u n g e t c _ n o l o c k . i n l                     _ u n g e t c _ n o l o c k         f:\dd\vctools\crt\crtw32\stdio\_file.c          (�<�L�    W a r n i n g       E r r o r       A s s e r t i o n   F a i l e d         . . .       m o d e   = =   _ C R T _ R P T H O O K _ I N S T A L L   | |   m o d e   = =   _ C R T _ R P T H O O K _ R E M O V E                           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ d b g r p t . c                     _ C r t S e t R e p o r t H o o k W 2           p f n N e w H o o k   ! =   N U L L             ( " T h e   h o o k   f u n c t i o n   i s   n o t   i n   t h e   l i s t ! " , 0 )                       f:\dd\vctools\crt\crtw32\misc\dbgrpt.c          _ _ c r t M e s s a g e W i n d o w W               w c s c p y _ s ( s z E x e N a m e ,   2 6 0 ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                       < p r o g r a m   n a m e   u n k n o w n >                 m e m c p y _ s ( s z S h o r t P r o g N a m e ,   s i z e o f ( T C H A R )   *   ( 2 6 0   -   ( s z S h o r t P r o g N a m e   -   s z E x e N a m e ) ) ,   d o t d o t d o t ,   s i z e o f ( T C H A R )   *   3 )                                                     
 
 F o r   i n f o r m a t i o n   o n   h o w   y o u r   p r o g r a m   c a n   c a u s e   a n   a s s e r t i o n 
 f a i l u r e ,   s e e   t h e   V i s u a l   C + +   d o c u m e n t a t i o n   o n   a s s e r t s .                                                 E x p r e s s i o n :           
 
     
 L i n e :         
 F i l e :         
 M o d u l e :             D e b u g   % s ! 
 
 P r o g r a m :   % s % s % s % s % s % s % s % s % s % s % s % s 
 
 ( P r e s s   R e t r y   t o   d e b u g   t h e   a p p l i c a t i o n ) 
                                       ( * _ e r r n o ( ) )           w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r                     M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y                 h�p�x�|���    Free    Normal  CRT Ignore  Client  _ C r t C h e c k M e m o r y ( )           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ d b g h e a p . c                   Client hook allocation failure at file %hs line %d.
            Client hook allocation failure.
        Invalid allocation size: %Iu bytes.
        Error: memory allocation: bad memory block type.
           Client hook re-allocation failure at file %hs line %d.
             Client hook re-allocation failure.
         Invalid allocation size: %Iu bytes.

Memory allocated at %hs(%d).
              Error: memory allocation: bad memory block type.

Memory allocated at %hs(%d).
                 The Block at 0x%p was allocated by aligned routines, use _aligned_realloc()                     _ C r t I s V a l i d H e a p P o i n t e r ( p U s e r D a t a )                       p O l d B l o c k - > n L i n e   = =   I G N O R E _ L I N E   & &   p O l d B l o c k - > l R e q u e s t   = =   I G N O R E _ R E Q                                 Error: possible heap corruption at or near 0x%p                 f R e a l l o c   | |   ( ! f R e a l l o c   & &   p N e w B l o c k   = =   p O l d B l o c k )                       _ p L a s t B l o c k   = =   p O l d B l o c k             _ p F i r s t B l o c k   = =   p O l d B l o c k               p U s e r D a t a   ! =   N U L L           _ e x p a n d _ d b g           The Block at 0x%p was allocated by aligned routines, use _aligned_free()                Client hook free failure.
      _ B L O C K _ T Y P E _ I S _ V A L I D ( p H e a d - > n B l o c k U s e )                     HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.

Memory allocated at %hs(%d).
                                         HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.
                               HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.

Memory allocated at %hs(%d).
                                     HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.
                           p H e a d - > n L i n e   = =   I G N O R E _ L I N E   & &   p H e a d - > l R e q u e s t   = =   I G N O R E _ R E Q                             p H e a d - > n B l o c k U s e   = =   n B l o c k U s e               _ p L a s t B l o c k   = =   p H e a d             _ p F i r s t B l o c k   = =   p H e a d           _ m s i z e _ d b g         _heapchk fails with _HEAPBADBEGIN.
         _heapchk fails with _HEAPBADNODE.
          _heapchk fails with _HEAPBADEND.
       _heapchk fails with _HEAPBADPTR.
       _heapchk fails with unknown return value!
          DAMAGED     HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.

Memory allocated at %hs(%d).
                                 HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.
                               %hs located at 0x%p is %Iu bytes long.

Memory allocated at %hs(%d).
               %hs located at 0x%p is %Iu bytes long.
             ( f N e w B i t s = = _ C R T D B G _ R E P O R T _ F L A G )   | |   ( ( f N e w B i t s   &   0 x 0 f f f f   &   ~ ( _ C R T D B G _ A L L O C _ M E M _ D F   |   _ C R T D B G _ D E L A Y _ F R E E _ M E M _ D F   |   _ C R T D B G _ C H E C K _ A L W A Y S _ D F   |   _ C R T D B G _ C H E C K _ C R T _ D F   |   _ C R T D B G _ L E A K _ C H E C K _ D F )   )   = =   0 )                                                                                 _ C r t S e t D b g F l a g         p f n   ! =   N U L L       _ C r t D o F o r A l l C l i e n t O b j e c t s               s t a t e   ! =   N U L L           _ C r t M e m C h e c k p o i n t           Bad memory block found at 0x%p.

Memory allocated at %hs(%d).
              Bad memory block found at 0x%p.
        _ C r t M e m D i f f e r e n c e           o l d S t a t e   ! =   N U L L         n e w S t a t e   ! =   N U L L         %.2X    _ p r i n t M e m B l o c k D a t a              Data: <%s> %s
     Dumping objects ->
     #File Error#(%d) :      %hs(%d) :       {%ld}   client block at 0x%p, subtype %x, %Iu bytes long.
              normal block at 0x%p, %Iu bytes long.
          crt block at 0x%p, subtype %x, %Iu bytes long.
             Object dump complete.
      Detected memory leaks!
     _ C r t M e m D u m p S t a t i s t i c s           %Id bytes in %Id %hs Blocks.
       Largest number used: %Id bytes.
        Total allocations: %Id bytes.
          I S _ 2 _ P O W _ N ( a l i g n )           _ a l i g n e d _ o f f s e t _ m a l l o c _ d b g             o f f s e t   = =   0   | |   o f f s e t   <   s i z e                 The block at 0x%p was not allocated by _aligned routines, use realloc()                 Damage before 0x%p which was allocated by aligned routine
              _ a l i g n e d _ o f f s e t _ r e a l l o c _ d b g                   The block at 0x%p was not allocated by _aligned routines, use free()                m e m b l o c k   ! =   N U L L         _ a l i g n e d _ m s i z e _ d b g             csm�               �                \@
R    �S    f:\dd\vctools\crt\crtw32\startup\dllcrt0.c                                    �A������               �             ��      �C      �C   ����G   ���8      `E           � 3  ?     �  ?                          f:\dd\vctools\crt\crtw32\startup\mlock.c            +;�@6X"l    bad exception                                                                                                                                                                                                                                                                                         ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               ( ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                                                            �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ w c s d u p . c                     _ w c s d u p _ d b g       w c s c p y _ s ( m e m o r y ,   s i z e ,   s t r i n g )                 f:\dd\vctools\crt\crtw32\misc\initctyp.c            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ i n i t c t y p . c                     p l o c i - > c t y p e 1 _ r e f c o u n t   >   0                 ( " C o r r u p t e d   p o i n t e r   p a s s e d   t o   _ f r e e a " ,   0 )                       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ m a l l o c . h                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ s e t l o c a l . c                     s e t l o c a l e           m b s t o w c s _ s ( & s i z e ,   ( ( v o i d   * ) 0 ) ,   0 ,   _ l o c a l e ,   2 1 4 7 4 8 3 6 4 7 )                         f:\dd\vctools\crt\crtw32\misc\setlocal.c            m b s t o w c s _ s ( ( ( v o i d   * ) 0 ) ,   i n w l o c a l e ,   s i z e ,   _ l o c a l e ,   ( ( s i z e _ t ) - 1 ) )                                   _ w c s t o m b s _ s _ l ( & s i z e ,   ( ( v o i d   * ) 0 ) ,   0 ,   o u t w l o c a l e ,   0 ,   & l o c a l e )                                 _ w c s t o m b s _ s _ l ( ( ( v o i d   * ) 0 ) ,   o u t l o c a l e ,   s i z e ,   o u t w l o c a l e ,   ( ( s i z e _ t ) - 1 ) ,   & l o c a l e )                                     ( ( p t l o c i - > l c _ c a t e g o r y [ _ c a t e g o r y ] . l o c a l e   ! =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ _ c a t e g o r y ] . r e f c o u n t   ! =   N U L L ) )   | |   ( ( p t l o c i - > l c _ c a t e g o r y [ _ c a t e g o r y ] . l o c a l e   = =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ _ c a t e g o r y ] . r e f c o u n t   = =   N U L L ) )                                                                                         ( f i l e   ! =   N U L L )             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f o p e n . c                     _ f s o p e n       ( m o d e   ! =   N U L L )         ( * m o d e   ! =   _ T ( ' \ 0 ' ) )           ( p f i l e   ! =   N U L L )           f o p e n _ s           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f s e e k . c                     f s e e k       _ w f s o p e n         _ w f o p e n _ s       k e r n e l 3 2 . d l l         FlsAlloc    FlsFree     FlsGetValue     FlsSetValue     InitializeCriticalSectionEx         CreateEventExW      CreateSemaphoreExW      SetThreadStackGuarantee     CreateThreadpoolTimer       SetThreadpoolTimer      WaitForThreadpoolTimerCallbacks         CloseThreadpoolTimer        CreateThreadpoolWait        SetThreadpoolWait       CloseThreadpoolWait     FlushProcessWriteBuffers        FreeLibraryWhenCallbackReturns          GetCurrentProcessorNumber       GetLogicalProcessorInformation          CreateSymbolicLinkW     SetDefaultDllDirectories        EnumSystemLocalesEx     CompareStringEx     GetDateFormatEx     GetLocaleInfoEx     GetTimeFormatEx     GetUserDefaultLocaleName        IsValidLocaleName       LCMapStringEx   GetCurrentPackageId     GetTickCount64      GetFileInformationByHandleExW       SetFileInformationByHandleW         ( f o r m a t   ! =   N U L L )             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ s p r i n t f . c                     s p r i n t f       ( s t r i n g   ! =   N U L L )         p V a l u e   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ d o s \ d o s m a p . c                   _ g e t _ e r r n o         _ g e t _ d o s e r r n o           f:\dd\vctools\crt\crtw32\time\strftime.c            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ t i m e \ s t r f t i m e . c                     _ G e t d a y s _ l         s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > w d a y _ a b b r [ n ] )                             s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > w d a y [ n ] )                       _ G e t m o n t h s _ l         s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > m o n t h _ a b b r [ n ] )                           s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > m o n t h [ n ] )                     (   s t r i n g   ! =   N U L L   )             _ S t r f t i m e _ l       (   m a x s i z e   ! =   0   )         (   f o r m a t   ! =   N U L L   )             (   t i m e p t r   ! =   N U L L   )           f:\dd\vctools\crt\crtw32\time\wcsftime.c            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ t i m e \ w c s f t i m e . c                     _ W _ G e t d a y s _ l             w c s c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > _ W _ w d a y _ a b b r [ n ] )                               w c s c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > _ W _ w d a y [ n ] )                         _ W _ G e t m o n t h s _ l             w c s c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > _ W _ m o n t h _ a b b r [ n ] )                             w c s c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > _ W _ m o n t h [ n ] )                       _ W _ G e t t n a m e s _ l             s t r c p y _ s ( d e s t - > w d a y _ a b b r [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > w d a y _ a b b r [ i d x ] )                                       s t r c p y _ s ( d e s t - > w d a y [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > w d a y [ i d x ] )                                   s t r c p y _ s ( d e s t - > m o n t h _ a b b r [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > m o n t h _ a b b r [ i d x ] )                                           s t r c p y _ s ( d e s t - > m o n t h [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > m o n t h [ i d x ] )                                       s t r c p y _ s ( d e s t - > a m p m [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > a m p m [ i d x ] )                                   s t r c p y _ s ( d e s t - > w w _ s d a t e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > w w _ s d a t e f m t )                                           s t r c p y _ s ( d e s t - > w w _ l d a t e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > w w _ l d a t e f m t )                                           s t r c p y _ s ( d e s t - > w w _ t i m e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > w w _ t i m e f m t )                                       w c s c p y _ s ( d e s t - > _ W _ w d a y _ a b b r [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w d a y _ a b b r [ i d x ] )                                             w c s c p y _ s ( d e s t - > _ W _ w d a y [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w d a y [ i d x ] )                                         w c s c p y _ s ( d e s t - > _ W _ m o n t h _ a b b r [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ m o n t h _ a b b r [ i d x ] )                                                 w c s c p y _ s ( d e s t - > _ W _ m o n t h [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ m o n t h [ i d x ] )                                             w c s c p y _ s ( d e s t - > _ W _ a m p m [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ a m p m [ i d x ] )                                         w c s c p y _ s ( d e s t - > _ W _ w w _ s d a t e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w w _ s d a t e f m t )                                         w c s c p y _ s ( d e s t - > _ W _ w w _ l d a t e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w w _ l d a t e f m t )                                         w c s c p y _ s ( d e s t - > _ W _ w w _ t i m e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w w _ t i m e f m t )                                             w c s c p y _ s ( d e s t - > _ W _ w w _ l o c a l e _ n a m e ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w w _ l o c a l e _ n a m e )                                             _ W c s f t i m e _ l       t i m e p t r   ! =   N U L L           F A L S E           (   (   t i m e p t r - > t m _ w d a y   > = 0   )   & &   (   t i m e p t r - > t m _ w d a y   < =   6   )   )                           _ W _ e x p a n d t i m e           (   (   t i m e p t r - > t m _ m o n   > = 0   )   & &   (   t i m e p t r - > t m _ m o n   < =   1 1   )   )                         (   (   t i m e p t r - > t m _ m d a y   > = 1   )   & &   (   t i m e p t r - > t m _ m d a y   < =   3 1   )   )                             (   (   t i m e p t r - > t m _ h o u r   > = 0   )   & &   (   t i m e p t r - > t m _ h o u r   < =   2 3   )   )                             (   (   t i m e p t r - > t m _ y d a y   > = 0   )   & &   (   t i m e p t r - > t m _ y d a y   < =   3 6 5   )   )                           (   (   t i m e p t r - > t m _ m i n   > = 0   )   & &   (   t i m e p t r - > t m _ m i n   < =   5 9   )   )                         (   (   t i m e p t r - > t m _ s e c   > = 0   )   & &   (   t i m e p t r - > t m _ s e c   < =   5 9   )   )                         (   t i m e p t r - > t m _ y e a r   > = 0   )                 (   t i m e p t r - > t m _ y e a r   > =   - 1 9 0 0   )   & &   (   t i m e p t r - > t m _ y e a r   < =   8 0 9 9   )                               _ m b s t o w c s _ s _ l ( & w n u m ,   * s t r i n g ,   * l e f t ,   ( _ _ t z n a m e ( ) ) [ ( ( t i m e p t r - > t m _ i s d s t ) ? 1 : 0 ) ] ,   ( ( s i z e _ t ) - 1 ) ,   p l o c i n f o )                                               (   " I n v a l i d   f o r m a t   d i r e c t i v e "   ,   0   )                 a m / p m       a / p       c c h C o u n t 1 = = 0   & &   c c h C o u n t 2 = = 1   | |   c c h C o u n t 1 = = 1   & &   c c h C o u n t 2 = = 0                                 f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ a _ c m p . c                   c a     z h - C H S     c s     d a     d e     e l     e n     e s     f i     f r     h e     h u     i s     i t     j a     k o     n l     n o     p l     p t     r o     r u     h r     s k     s q     s v     t h     t r     u r     i d     u k     b e     s l     e t     l v     l t     f a     v i     h y     a z     e u     m k     a f     k a     f o     h i     m s     k k     k y     s w     u z     t t     p a     g u     t a     t e     k n     m r     s a     m n     g l     k o k       s y r       d i v       a r - S A       b g - B G       c a - E S       z h - T W       c s - C Z       d a - D K       d e - D E       e l - G R       e n - U S       f i - F I       f r - F R       h e - I L       h u - H U       i s - I S       i t - I T       j a - J P       k o - K R       n l - N L       n b - N O       p l - P L       p t - B R       r o - R O       r u - R U       h r - H R       s k - S K       s q - A L       s v - S E       t h - T H       t r - T R       u r - P K       i d - I D       u k - U A       b e - B Y       s l - S I       e t - E E       l v - L V       l t - L T       f a - I R       v i - V N       h y - A M       a z - A Z - L a t n         e u - E S       m k - M K       t n - Z A       x h - Z A       z u - Z A       a f - Z A       k a - G E       f o - F O       h i - I N       m t - M T       s e - N O       m s - M Y       k k - K Z       k y - K G       s w - K E       u z - U Z - L a t n         t t - R U       b n - I N       p a - I N       g u - I N       t a - I N       t e - I N       k n - I N       m l - I N       m r - I N       s a - I N       m n - M N       c y - G B       g l - E S       k o k - I N     s y r - S Y     d i v - M V     q u z - B O     n s - Z A       m i - N Z       a r - I Q       z h - C N       d e - C H       e n - G B       e s - M X       f r - B E       i t - C H       n l - B E       n n - N O       p t - P T       s r - S P - L a t n         s v - F I       a z - A Z - C y r l         s e - S E       m s - B N       u z - U Z - C y r l         q u z - E C     a r - E G       z h - H K       d e - A T       e n - A U       e s - E S       f r - C A       s r - S P - C y r l         s e - F I       q u z - P E     a r - L Y       z h - S G       d e - L U       e n - C A       e s - G T       f r - C H       h r - B A       s m j - N O     a r - D Z       z h - M O       d e - L I       e n - N Z       e s - C R       f r - L U       b s - B A - L a t n         s m j - S E     a r - M A       e n - I E       e s - P A       f r - M C       s r - B A - L a t n         s m a - N O     a r - T N       e n - Z A       e s - D O       s r - B A - C y r l         s m a - S E     a r - O M       e n - J M       e s - V E       s m s - F I     a r - Y E       e n - C B       e s - C O       s m n - F I     a r - S Y       e n - B Z       e s - P E       a r - J O       e n - T T       e s - A R       a r - L B       e n - Z W       e s - E C       a r - K W       e n - P H       e s - C L       a r - A E       e s - U Y       a r - B H       e s - P Y       a r - Q A       e s - B O       e s - S V       e s - H N       e s - N I       e s - P R       z h - C H T     s r         p�B   $,   t5q   �?    �5�   �5�   �5�   �5�   �5�   �5�   �5�   �5�   6�   6�   $6�   46�   D6C   T6�   d6�   t6�   )   �6�   �6k   �!   �6c   �?   �6D   �6}   �6�   �   7E   �   7G   (7�   �   87H   �   H7�   X7�   h7I   x7�   �7�   �A   �7�   �   �7J      �7�   �7�   �7�   �7�   �7�   8�   8�   (8�   88�   H8�   X8K   h8�   x8�   	   �8�   �8�   �8�   �8�   �8�   �8�   �8�   �8�   9�   9�   (9�   89�   H9�   X9�   h9�   x9�   �9�   �9�   �9�   �#   �9e   *   �9l   �&   �9h   
   �9L   4.   �9s      :�   :�   (:�   8:M   H:�   X:�   �>   h:�   |7   x:   $   �:N   </   �:t   �   �:�   �:Z   ,   �:O   (   �:j   �   �:a   4   �:P   <   ;�   ;Q   D   (;R   ,-   8;r   L1   H;x   �:   X;�   L   �?   h;�   x;S   T2   �;y   �%   �;g   �$   �;f   �;�   +   �;m   �;�   �=   �;�   �;   �;�   D0   <�   <w   (<u   8<U   T   H<�   X<T   h<�   \   x<�   t6   �<~   d   �<V   l   �<W   �<�   �<�   �<�   �<�   t   �<X   |   =Y   �<   =�   (=�   8=v   H=�   �   X=[   �"   h=d   x=�   �=�   �=�   �=�   �=�   �=�   �   �=\   L$�   �=�   >�    >�   <>�   �   X>�   h>]   \3   x>z   �@   �>�   �8   �>�   �9   �>�   �   �>^   �>n   �   �>_   l5   �>|   �    �>b   �   ?`   d4   ?�   4?{   �'   P?i   `?o   p?   �?�   �?�   �?�   �?�   �?�   �?F   �?p      �?   �?   �   �   �   �   �   �	   
            $   ,   4   <   D   L   T   \   d   l   t   |   �   �   �   �   �   �    �!   �"   �#   �$   �%   �&   �'   �)   �*   �+   ,   -   /   6   $7   ,8   49   <>   D?   L@   TA   \C   dD   lF   tG   |I   �J   �K   �N   �O   �P   �V   �W   �Z   �e   �   p�  �  �          0  @  P	  `  p  �  �  �  �  �  �  �  �          0  @  P  `  p  �  �  �   �!  �"  �#  �$  �%   &  '   )  0*  @+  P,  `-  |/  �2  �4  �5  �6  �7  �8  �9  �:  ;  >  ,?  <@  LA  \C  lD  �E  �F  �G  �I  �J  �K  �L  �N  O  P  (R  8V  HW  XZ  he  xk  �l  ��  �  �  �  �	  �
  �      (  8  H  X  t,  �;  �>  �C  �k  �  �  �   	   
  ,   <   L ;  h k  x   �   �   � 	  � 
  �   �   � ;  �   !  !  (!	  8!
  H!  X!  h!;  �!  �!	  �!
  �!  �!  �!;  �!   "	  "
   "  0";  L"   \"	   l"
   |";   �"$  �"	$  �"
$  �";$  �"(  �"	(  �"
(  �",  #	,  #
,  ,#0  <#	0  L#
0  \#4  l#	4  |#
4  �#8  �#
8  �#<  �#
<  �#@  �#
@  �#
D  �#
H  $
L  $
P  ,$|  <$|  L$                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            a f - z a       a r - a e       a r - b h       a r - d z       a r - e g       a r - i q       a r - j o       a r - k w       a r - l b       a r - l y       a r - m a       a r - o m       a r - q a       a r - s a       a r - s y       a r - t n       a r - y e       a z - a z - c y r l         a z - a z - l a t n         b e - b y       b g - b g       b n - i n       b s - b a - l a t n         c a - e s       c s - c z       c y - g b       d a - d k       d e - a t       d e - c h       d e - d e       d e - l i       d e - l u       d i v - m v     e l - g r       e n - a u       e n - b z       e n - c a       e n - c b       e n - g b       e n - i e       e n - j m       e n - n z       e n - p h       e n - t t       e n - u s       e n - z a       e n - z w       e s - a r       e s - b o       e s - c l       e s - c o       e s - c r       e s - d o       e s - e c       e s - e s       e s - g t       e s - h n       e s - m x       e s - n i       e s - p a       e s - p e       e s - p r       e s - p y       e s - s v       e s - u y       e s - v e       e t - e e       e u - e s       f a - i r       f i - f i       f o - f o       f r - b e       f r - c a       f r - c h       f r - f r       f r - l u       f r - m c       g l - e s       g u - i n       h e - i l       h i - i n       h r - b a       h r - h r       h u - h u       h y - a m       i d - i d       i s - i s       i t - c h       i t - i t       j a - j p       k a - g e       k k - k z       k n - i n       k o k - i n     k o - k r       k y - k g       l t - l t       l v - l v       m i - n z       m k - m k       m l - i n       m n - m n       m r - i n       m s - b n       m s - m y       m t - m t       n b - n o       n l - b e       n l - n l       n n - n o       n s - z a       p a - i n       p l - p l       p t - b r       p t - p t       q u z - b o     q u z - e c     q u z - p e     r o - r o       r u - r u       s a - i n       s e - f i       s e - n o       s e - s e       s k - s k       s l - s i       s m a - n o     s m a - s e     s m j - n o     s m j - s e     s m n - f i     s m s - f i     s q - a l       s r - b a - c y r l         s r - b a - l a t n         s r - s p - c y r l         s r - s p - l a t n         s v - f i       s v - s e       s w - k e       s y r - s y     t a - i n       t e - i n       t h - t h       t n - z a       t r - t r       t t - r u       u k - u a       u r - p k       u z - u z - c y r l         u z - u z - l a t n         v i - v n       x h - z a       z h - c h s     z h - c h t     z h - c n       z h - h k       z h - m o       z h - s g       z h - t w       z u - z a       a r     b g     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ w i n a p i n l s . c                   _ _ c r t D o w n l e v e l L C I D T o L o c a l e N a m e                 w c s c p y _ s ( o u t L o c a l e N a m e ,   c c h L o c a l e N a m e ,   b u f f e r )                     �A�BHDlD�D�D                   Stack around the variable ' ' was corrupted.    The variable '  ' is being used without being initialized.                                      The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.
                                                    A cast to a smaller data type has caused a loss of data.  If this was intentional, you should mask the source of the cast with the appropriate bitmask.  For example:  
	char c = (i & 0xFF);
Changing the code in this way will not affect the quality of the resulting optimized code.
                                                            Stack memory was corrupted
        A local variable was used before it was initialized
           Stack memory around _alloca was corrupted
         Unknown Runtime Check Error
           R u n t i m e   C h e c k   E r r o r . 
    U n a b l e   t o   d i s p l a y   R T C   M e s s a g e .                               R u n - T i m e   C h e c k   F a i l u r e   # % d   -   % s               Unknown Filename    Unknown Module Name     Run-Time Check Failure #%d - %s         Stack corrupted near unknown variable           u s e r 3 2 . d l l         wsprintfA   Stack area around _alloca memory reserved by this function is corrupted
                
Data: <    
Allocation number within this function:            
Size:      
Address: 0x        Stack area around _alloca memory reserved by this function is corrupted                 %s%s%p%s%ld%s%d%s       
   >   %s%s%s%s    A variable is being used without being initialized.             H<HpH�H�H    Stack pointer corruption        Cast to smaller type causing loss of data           Stack memory corruption     Local variable used before initialization           Stack around _alloca corrupted          The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.                                              f:\dd\vctools\crt\crtw32\misc\i386\chkesp.c                K   xK	   �K
   PL   �L   M   �M   �M   @N   �N    O   �O    P   xP   �P    �Q!   8R"   �Tx   Uy   (Uz   HU�   lU�   tU                                        R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
                         R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
                       R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
                           R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
                     R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
                           R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
                         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
                 R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
                         R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
                         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
                       R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
                         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
                         R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
                 R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
                     R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
                                             R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
                             R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
                                                                                                     R 6 0 3 4  
 -   i n c o n s i s t e n t   o n e x i t   b e g i n - e n d   v a r i a b l e s  
                         D O M A I N   e r r o r  
         S I N G   e r r o r  
         T L O S S   e r r o r  
            
     r u n t i m e   e r r o r           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t a r t u p \ c r t 0 m s g . c                     _ N M S G _ W R I T E           w c s c p y _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " R u n t i m e   E r r o r ! \ n \ n P r o g r a m :   " )                                     R u n t i m e   E r r o r ! 
 
 P r o g r a m :                 w c s c p y _ s ( p r o g n a m e ,   p r o g n a m e _ s i z e ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                                 w c s n c p y _ s ( p c h ,   p r o g n a m e _ s i z e   -   ( p c h   -   p r o g n a m e ) ,   L " . . . " ,   3 )                           w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " \ n \ n " )                                   w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   e r r o r _ t e x t )                             f:\dd\vctools\crt\crtw32\misc\inithelp.c                f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ i n i t h e l p . c                     _ _ g e t l o c a l e i n f o               s t r n c p y _ s ( * s t r a d d r e s s ,   o u t s i z e ,   p c b u f f e r ,   o u t s i z e   -   1 )                         m s c o r e e . d l l       CorExitProcess          f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t a r t u p \ c r t 0 d a t . c                     _ g e t _ w p g m p t r         _ w p g m p t r   ! =   N U L L         _ g e t _ p g m p t r       _ p g m p t r   ! =   N U L L           p a t h   ! =   N U L L         _ _ c o p y _ p a t h _ t o _ w i d e _ s t r i n g             o u t P a t h   ! =   N U L L           f:\dd\vctools\crt\crtw32\startup\crt0dat.c          i n S t r i n g   ! =   N U L L         _ _ c o p y _ t o _ c h a r         o u t S t r i n g   ! =   N U L L           exp pow log log10   sinh    cosh    tanh    asin    acos    atan    atan2   sqrt    sin cos tan ceil    floor   fabs    modf    ldexp   _cabs   _hypot  fmod    frexp   _y0 _y1 _yn _logb   _nextafter          ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n B y t e s ) )   >   0                         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ t c s c p y _ s . i n l                   s t r c p y _ s         ( ( ( _ S r c ) ) )   ! =   N U L L             B u f f e r   i s   t o o   s m a l l           ( L " B u f f e r   i s   t o o   s m a l l "   & &   0 )               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f i l e n o . c                   _ f i l e n o           ( f h   > =   0   & &   ( u n s i g n e d ) f h   <   ( u n s i g n e d ) _ n h a n d l e )                     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ c l o s e . c                     _ c l o s e     ( _ o s f i l e ( f h )   &   F O P E N )               ( " I n v a l i d   f i l e   d e s c r i p t o r .   F i l e   p o s s i b l y   c l o s e d   b y   a   d i f f e r e n t   t h r e a d " , 0 )                                   s t r e a m   ! =   N U L L         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ f r e e b u f . c                       ( f i l e d e s   > =   0   & &   ( u n s i g n e d ) f i l e d e s   <   ( u n s i g n e d ) _ n h a n d l e )                         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ c o m m i t . c                   _ c o m m i t       ( _ o s f i l e ( f i l e d e s )   &   F O P E N )                 f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ w r i t e . c                     _ w r i t e     ( b u f   ! =   N U L L )           _ w r i t e _ n o l o c k           ( ( c n t   &   1 )   = =   0 )         i s l e a d b y t e ( _ d b c s B u f f e r ( f h ) )                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ f i l b u f . c                     _ f i l b u f       f:\dd\vctools\crt\crtw32\lowio\ioinit.c         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f t e l l i 6 4 . c                   _ f t e l l i 6 4           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ f l s b u f . c                         ( " i n c o n s i s t e n t   I O B   f i e l d s " ,   s t r e a m - > _ p t r   -   s t r e a m - > _ b a s e   > =   0 )                             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ l s e e k i 6 4 . c                   _ l s e e k i 6 4           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ g e t b u f . c                     f:\dd\vctools\crt\crtw32\stdio\_getbuf.c            ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n W o r d s ) )   >   0                     w c s c p y _ s             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ s w p r i n t f . c                   _ s w p r i n t f       f:\dd\vctools\crt\crtw32\misc\winsig.c          ( " I n v a l i d   s i g n a l   o r   e r r o r " ,   0 )                 f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ w i n s i g . c                     s i g n a l     r a i s e       U S E R 3 2 . D L L         MessageBoxW     GetActiveWindow     GetLastActivePopup      GetUserObjectInformationW       GetProcessWindowStation         n R p t T y p e   > =   0   & &   n R p t T y p e   <   _ C R T _ E R R C N T                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ d b g r p t t . c                   _ C r t S e t R e p o r t M o d e               f M o d e   = =   _ C R T D B G _ R E P O R T _ M O D E   | |   ( f M o d e   &   ~ ( _ C R T D B G _ M O D E _ F I L E   |   _ C R T D B G _ M O D E _ D E B U G   |   _ C R T D B G _ M O D E _ W N D W ) )   = =   0                                                 _ C r t S e t R e p o r t F i l e           _ V C r t D b g R e p o r t A               _ i t o a _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   Second Chance Assertion Failed: File            <file unknown>      , Line      s t r c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   _CrtDbgReport: String too long or IO Error              s t r c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   " A s s e r t i o n   f a i l e d :   "   :   " A s s e r t i o n   f a i l e d ! " )                                     Assertion failed:       Assertion failed!           s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ r " )                          s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ n " )                   %s(%d) : %s     s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                     s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                           e   =   m b s t o w c s _ s ( & r e t ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               w c s c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                         _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g                             _ V C r t D b g R e p o r t W           _ i t o w _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   S e c o n d   C h a n c e   A s s e r t i o n   F a i l e d :   F i l e                     < f i l e   u n k n o w n >         ,   L i n e         
   w c s c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                 w c s c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   L " A s s e r t i o n   f a i l e d :   "   :   L " A s s e r t i o n   f a i l e d ! " )                                     A s s e r t i o n   f a i l e d :               A s s e r t i o n   f a i l e d !               w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ r " )                        w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ n " )                 % s ( % d )   :   % s           w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                           w c s t o m b s _ s ( ( ( v o i d   * ) 0 ) ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                                 s t r c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                           _CrtDbgReport: String too long or Invalid characters in String                  w c s t o m b s _ s ( & r e t ,   s z a O u t M e s s a g e ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . l o c a l e   ! =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . r e f c o u n t   ! =   N U L L ) )   | |   ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . l o c a l e   = =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . r e f c o u n t   = =   N U L L ) )                                                                                         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ l o c a l r e f . c                     ���    f:\dd\vctools\crt\crtw32\mbstring\mbctype.c         c   > =   - 1   & &   c   < =   2 5 5               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ i s c t y p e . c                     p B l o c k   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h e a p \ e x p a n d . c                     _ e x p a n d _ b a s e         (�<�L�    ... _ C r t S e t R e p o r t H o o k 2             _ _ c r t M e s s a g e W i n d o w A               s t r c p y _ s ( s z E x e N a m e ,   2 6 0 ,   " < p r o g r a m   n a m e   u n k n o w n > " )                         <program name unknown>      D e b u g   % s ! 
 
 P r o g r a m :   % h s % s % s % h s % s % h s % s % h s % s % s % h s % s 
 
 ( P r e s s   R e t r y   t o   d e b u g   t h e   a p p l i c a t i o n ) 
                                         f:\dd\vctools\crt\crtw32\startup\tidtable.c         p n h   = =   0         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h e a p \ h a n d l e r . c p p                   Sun Mon Tue Wed Thu Fri Sat Sunday  Monday  Tuesday     Wednesday   Thursday    Friday  Saturday    Jan Feb Mar Apr May Jun Jul Aug Sep Oct Nov Dec January     February    March   April   June    July    August  September   October     November    December    AM  PM  MM/dd/yy    dddd, MMMM dd, yyyy     HH:mm:ss    S u n       M o n       T u e       W e d       T h u       F r i       S a t       S u n d a y     M o n d a y     T u e s d a y       W e d n e s d a y       T h u r s d a y         F r i d a y     S a t u r d a y         J a n       F e b       M a r       A p r       M a y       J u n       J u l       A u g       S e p       O c t       N o v       D e c       J a n u a r y       F e b r u a r y         M a r c h       A p r i l       J u n e     J u l y     A u g u s t     S e p t e m b e r       O c t o b e r       N o v e m b e r         D e c e m b e r         A M     P M     M M / d d / y y         d d d d ,   M M M M   d d ,   y y y y           H H : m m : s s         _ c r t h e a p         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h e a p \ h e a p i n i t . c                     p N o d e - > _ N e x t   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ e h \ t y p n a m e . c p p                   t y p e _ i n f o : : _ N a m e _ b a s e               s t r c p y _ s   ( ( c h a r   * ) ( ( t y p e _ i n f o   * ) _ T h i s ) - > _ M _ d a t a ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                                 t y p e _ i n f o : : _ N a m e _ b a s e _ i n t e r n a l                     s t r c p y _ s   ( p T m p T y p e N a m e ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                       b u f   ! =   N U L L       f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ c o n v \ c v t . c                 _ c f t o e 2 _ l       s i z e I n B y t e s   >   0               s i z e I n B y t e s   >   ( s i z e _ t ) ( 3   +   ( n d e c   >   0   ?   n d e c   :   0 )   +   5   +   1 )                               s t r c p y _ s ( p ,   ( s i z e I n B y t e s   = =   ( s i z e _ t ) - 1   ?   s i z e I n B y t e s   :   s i z e I n B y t e s   -   ( p   -   b u f ) ) ,   " e + 0 0 0 " )                                       e+000   _ c f t o e _ l         _ c f t o a _ l         s i z e I n B y t e s   >   ( s i z e _ t ) ( 1   +   4   +   n d e c   +   6 )                     _ c f t o f 2 _ l       _ c f t o f _ l         _ c f t o g _ l             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t a r t u p \ i 3 8 6 \ f p 8 . c                       _ s e t d e f a u l t p r e c i s i o n             _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   0 x 0 0 0 1 0 0 0 0 ,   0 x 0 0 0 3 0 0 0 0 )                         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          �      	                                   f:\dd\vctools\crt\crtw32\startup\stdargv.c          f:\dd\vctools\crt\crtw32\startup\stdenvp.c          f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t a r t u p \ s t d e n v p . c                     _ s e t e n v p         s t r c p y _ s ( * e n v ,   c c h a r s ,   p )               f:\dd\vctools\crt\crtw32\misc\a_env.c           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ v s p r i n t f . c                   _ v s n p r i n t f _ l             ( c o u n t   = =   0 )   | |   ( s t r i n g   ! =   N U L L )                        ���5�h!����?      �?                            �?5�h!���>@�������             ��      �@      �                            ��    �H�����E�����MԐ��.����\����'                L C _ A L L     L C _ C O L L A T E         L C _ C T Y P E         L C _ M O N E T A R Y       L C _ N U M E R I C         L C _ T I M E       	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~                         ( " I n v a l i d   p a r a m e t e r   f o r   _ c o n f i g t h r e a d l o c a l e " , 0 )                           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ w s e t l o c a . c                     _ c o n f i g t h r e a d l o c a l e           f:\dd\vctools\crt\crtw32\misc\wsetloca.c            L C _ M I N   < =   _ c a t e g o r y   & &   _ c a t e g o r y   < =   L C _ M A X                     _ w s e t l o c a l e       = ;     ;   _ w s e t l o c a l e _ n o l o c k             w c s n c p y _ s ( l c t e m p ,   ( s i z e o f ( l c t e m p )   /   s i z e o f ( l c t e m p [ 0 ] ) ) ,   s ,   l e n )                               _ w s e t l o c a l e _ s e t _ c a t               w c s c p y _ s ( p c h _ c a t _ l o c a l e ,   c c h ,   l c t e m p )                   =   _ w s e t l o c a l e _ g e t _ a l l           w c s c a t _ s ( p c h ,   c c h ,   L " ; " )             _ e x p a n d l o c a l e           w c s n c p y _ s ( l o c a l e N a m e O u t p u t ,   l o c a l e N a m e S i z e I n C h a r s , _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   ( s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   /   s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e [ 0 ] ) ) )                                                                             w c s c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   L " C " )                   C       w c s n c p y _ s ( l o c a l e N a m e O u t p u t ,   l o c a l e N a m e S i z e I n C h a r s ,   n a m e s . s z L o c a l e N a m e ,   w c s l e n ( n a m e s . s z L o c a l e N a m e )   +   1 )                                             w c s n c p y _ s ( c a c h e o u t ,   c a c h e o u t L e n ,   e x p r ,   c h a r a c t e r s I n E x p r e s s i o n   +   1 )                             w c s n c p y _ s ( l o c a l e N a m e O u t p u t ,   l o c a l e N a m e S i z e I n C h a r s ,   e x p r ,   c h a r a c t e r s I n E x p r e s s i o n   +   1 )                                         w c s n c p y _ s ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   ( s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   /   s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e [ 0 ] ) ) ,   e x p r ,   c h a r a c t e r s I n E x p r e s s i o n   +   1 )                                                                         w c s n c p y _ s ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   ( s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   /   s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e [ 0 ] ) ) ,   l o c a l e N a m e O u t p u t ,   w c s l e n ( l o c a l e N a m e O u t p u t )   +   1 )                                                                             w c s n c p y _ s ( c a c h e i n ,   c a c h e i n L e n ,   e x p r ,   c h a r a c t e r s I n E x p r e s s i o n   +   1 )                                 w c s c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   c a c h e o u t )                   _ w c s c a t s         w c s c a t _ s ( o u t s t r ,   n u m b e r O f E l e m e n t s ,   (   * ( w c h a r _ t   *   * ) ( ( s u b s t r   + =   (   ( s i z e o f ( w c h a r _ t   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   -   (   ( s i z e o f ( w c h a r _ t   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   ) )                                                                                   _ _ l c _ w c s t o l c         w c s n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   & w l o c a l e [ 1 ] ,   1 6 - 1 )                                               _ . ,       w c s n c p y _ s ( n a m e s - > s z L a n g u a g e ,   ( s i z e o f ( n a m e s - > s z L a n g u a g e )   /   s i z e o f ( n a m e s - > s z L a n g u a g e [ 0 ] ) ) ,   w l o c a l e ,   l e n )                                             w c s n c p y _ s ( n a m e s - > s z C o u n t r y ,   ( s i z e o f ( n a m e s - > s z C o u n t r y )   /   s i z e o f ( n a m e s - > s z C o u n t r y [ 0 ] ) ) ,   w l o c a l e ,   l e n )                                           w c s n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   w l o c a l e ,   l e n )                                             _ _ l c _ l c t o w c s         w c s c p y _ s ( l o c a l e ,   n u m b e r O f E l e m e n t s ,   n a m e s - > s z L a n g u a g e )                           _   .   _ _ c o p y _ l o c a l e _ n a m e                 w c s n c p y _ s ( l o c a l e N a m e C o p y ,   c c h + 1 ,   l o c a l e N a m e ,   c c h + 1 )                       s   ! =   N U L L           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ m b s t o w c s . c                       _ m b s t o w c s _ l _ h e l p e r                 ( p w c s   = =   N U L L   & &   s i z e I n W o r d s   = =   0 )   | |   ( p w c s   ! =   N U L L   & &   s i z e I n W o r d s   >   0 )                               _ m b s t o w c s _ s _ l           b u f f e r S i z e   < =   I N T _ M A X           r e t s i z e   < =   s i z e I n W o r d s             p w c s   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ w c s t o m b s . c                       _ w c s t o m b s _ l _ h e l p e r                 ( d s t   ! =   N U L L   & &   s i z e I n B y t e s   >   0 )   | |   ( d s t   = =   N U L L   & &   s i z e I n B y t e s   = =   0 )                               _ w c s t o m b s _ s _ l           s i z e I n B y t e s   >   r e t s i z e           f:\dd\vctools\crt\crtw32\stdio\stream.c         ccs UTF-8   UTF-16LE    UNICODE         f i l e n a m e   ! =   N U L L         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ o p e n . c                     m o d e   ! =   N U L L         ( " I n v a l i d   f i l e   o p e n   m o d e " , 0 )                 _ o p e n f i l e       ( * m o d e   = =   _ T ( ' \ 0 ' ) )           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f t e l l . c                     f t e l l       _ f t e l l _ n o l o c k               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ l s e e k . c                     _ l s e e k     ( " I n v a l i d   f i l e   d e s c r i p t o r " , 0 )               c c s   U T F - 8   U T F - 1 6 L E     U N I C O D E               _ w o p e n f i l e         _ v s p r i n t f _ l       _ v s c p r i n t f _ h e l p e r           _ v s n p r i n t f _ h e l p e r           f o r m a t   ! =   N U L L         _ v s p r i n t f _ s _ l               s t r i n g   ! =   N U L L   & &   s i z e I n B y t e s   >   0                   ( " B u f f e r   t o o   s m a l l " ,   0 )               _ v s n p r i n t f _ s _ l         (null)  ( n u l l )                EEE50 P    ( 8PX 700WP        `h````  xpxxxx                              f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ o u t p u t . c                   _ o u t p u t _ l       ( c h   ! =   _ T ( ' \ 0 ' ) )         ( " ' n '   f o r m a t   s p e c i f i e r   d i s a b l e d " ,   0 )                 f:\dd\vctools\crt\crtw32\stdio\output.c         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ w c s i c m p . c                   _ w c s i c m p _ l         _ w c s i c m p         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ t i m e \ t z s e t . c                   _ t z s e t _ n o l o c k           _ g e t _ t i m e z o n e ( & t i m e z o n e )             _ g e t _ d a y l i g h t ( & d a y l i g h t )             _ g e t _ d s t b i a s ( & d s t b i a s )             TZ  f:\dd\vctools\crt\crtw32\time\tzset.c               s t r c p y _ s ( l a s t T Z ,   s t r l e n ( T Z )   +   1 ,   T Z )                 s t r n c p y _ s ( t z n a m e [ 0 ] ,   6 4 ,   T Z ,   3 )                   s t r n c p y _ s ( t z n a m e [ 1 ] ,   6 4 ,   T Z ,   3 )               c v t d a t e       _ i s i n d s t _ n o l o c k           SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec                ( _ D a y l i g h t   ! =   N U L L )               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ t i m e \ t i m e s e t . c                   _ g e t _ d a y l i g h t               ( _ D a y l i g h t _ s a v i n g s _ b i a s   ! =   N U L L )                 _ g e t _ d s t b i a s         ( _ T i m e z o n e   ! =   N U L L )           _ g e t _ t i m e z o n e               ( _ B u f f e r   ! =   N U L L   & &   _ S i z e I n B y t e s   >   0 )   | |   ( _ B u f f e r   = =   N U L L   & &   _ S i z e I n B y t e s   = =   0 )                                   _ g e t _ t z n a m e       _ R e t u r n V a l u e   ! =   N U L L             _ I n d e x   = =   0   | |   _ I n d e x   = =   1             M S V C R 1 2 0 D . d l l   b i n \ M S P D B 1 2 0 . D L L                          ���   ��� �  A D V A P I 3 2 . D L L         RegOpenKeyExW   RegQueryValueExW    RegCloseKey         S O F T W A R E \ M i c r o s o f t \ V i s u a l S t u d i o \ 1 2 . 0 \ S e t u p \ V C                       P r o d u c t D i r         D L L       M S P D B 1 2 0         M S P D B 1 2 0         PDBOpenValidate5        f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ t c s c a t _ s . i n l                   w c s c a t _ s         S t r i n g   i s   n o t   n u l l   t e r m i n a t e d               ( L " S t r i n g   i s   n o t   n u l l   t e r m i n a t e d "   & &   0 )                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ t c s n c p y _ s . i n l                     w c s n c p y _ s       ( " I n v a l i d   e r r o r _ m o d e " ,   0 )                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ e r r m o d e . c                   _ s e t _ e r r o r _ m o d e           s t r n c p y _ s       _ R a n d o m V a l u e   ! =   N U L L                 f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ r a n d _ s . c                     r a n d _ s     ( " r a n d _ s   i s   n o t   a v a i l a b l e   o n   t h i s   p l a t f o r m " ,   0 )                       SystemFunction036           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ s f t b u f . c                     f:\dd\vctools\crt\crtw32\stdio\_sftbuf.c            f l a g   = =   0   | |   f l a g   = =   1             f:\dd\vctools\crt\crtw32\lowio\osfinfo.c                f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ o s f i n f o . c                     _ g e t _ o s f h a n d l e         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ i s a t t y . c                   _ i s a t t y           _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   1   | |   _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   2                                                 f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ m b t o w c . c                       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ r e a d . c                   _ r e a d       ( c n t   < =   I N T _ M A X )         _ r e a d _ n o l o c k         ( i n p u t b u f   ! =   N U L L )             f:\dd\vctools\crt\crtw32\lowio\read.c               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ v s w p r i n t . c                   _ v s w p r i n t f _ l         _ v s c w p r i n t f _ h e l p e r             _ v s w p r i n t f _ h e l p e r           _ v s w p r i n t f _ s _ l             s t r i n g   ! =   N U L L   & &   s i z e I n W o r d s   >   0                   _ v s n w p r i n t f _ s _ l           _ w o u t p u t _ l         s t r c a t _ s         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ x t o a . c                   x t o a _ s     s i z e I n T C h a r s   >   0         s i z e I n T C h a r s   >   ( s i z e _ t ) ( i s _ n e g   ?   2   :   1 )                   2   < =   r a d i x   & &   r a d i x   < =   3 6               l e n g t h   <   s i z e I n T C h a r s           x 6 4 t o a _ s         x t o w _ s     x 6 4 t o w _ s         f:\dd\vctools\crt\crtw32\misc\initmon.c         p l o c i - > l c o n v _ m o n _ r e f c o u n t   >   0                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ i n i t m o n . c                   f:\dd\vctools\crt\crtw32\misc\initnum.c         p l o c i - > l c o n v _ n u m _ r e f c o u n t   >   0               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ i n i t n u m . c                   f:\dd\vctools\crt\crtw32\misc\inittime.c                p l o c i - > l c _ t i m e _ c u r r - > r e f c o u n t   >   0                       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ i n i t t i m e . c                         ��������������(�0�<�L�\��ah�p�|����������������������������������������������������������������� �������$�0�<�H�d�p����������<�h��������(�<�@�H�\�������������$�P���������(�\����a�������,�                                                                                __based(    __cdecl     __pascal    __stdcall   __thiscall      __fastcall      __vectorcall    __clrcall   __eabi  __ptr64     __restrict      __unaligned     restrict(    new     delete     =   >>  <<  !   ==  !=  []  operator    ->  ++  --  +   &   ->* /   %   <   <=  >   >=  ,   ()  ~   ^   |   &&  ||  *=  +=  -=  /=  %=  >>= <<= &=  |=  ^=  `vftable'   `vbtable'   `vcall'     `typeof'    `local static guard'        `string'    `vbase destructor'      `vector deleting destructor'        `default constructor closure'       `scalar deleting destructor'        `vector constructor iterator'       `vector destructor iterator'        `vector vbase constructor iterator'         `virtual displacement map'      `eh vector constructor iterator'        `eh vector destructor iterator'         `eh vector vbase constructor iterator'          `copy constructor closure'      `udt returning'     `EH `RTTI   `local vftable'     `local vftable constructor closure'          new[]   delete[]   `omni callsig'      `placement delete closure'      `placement delete[] closure'        `managed vector constructor iterator'           `managed vector destructor iterator'        `eh vector copy constructor iterator'           `eh vector vbase copy constructor iterator'         `dynamic initializer for '      `dynamic atexit destructor for '        `vector copy constructor iterator'          `vector vbase copy constructor iterator'            `managed vector copy constructor iterator'          `local static thread guard'          Type Descriptor'        Base Class Descriptor at (          Base Class Array'       Class Hierarchy Descriptor'         Complete Object Locator'       CV:     ::  template-parameter-     generic-type-   `   '   `anonymous namespace'       ''  `non-type-template-parameter        void    `template-parameter     NULL    }'  }'  `vtordispex{    `vtordisp{      `adjustor{      `local static destructor helper'        `template static data member constructor helper'            `template static data member destructor helper'             static      virtual     private:    protected:      public:     [thunk]:    extern "C"      )   char    short   int     long    unsigned    void    volatile    std::nullptr_t      <ellipsis>      ,...    ,<ellipsis>      throw(     cpu amp ,   char    short   int long    float   double  bool    __int8  __int16     __int32     __int64     __int128    <unknown>   wchar_t     __w64   UNKNOWN     signed      const    volatile   `unknown ecsu'      union   struct      class   coclass     cointerface     enum    volatile    const   cli::array<     cli::pin_ptr<   )[  {flat}  {for    s   A�_�_�_    hA�j%n&6    �Al`B@     B�Y�>�j    |BG[�Ms    �B�\�N�=     ??     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ _ f p t o s t r . c                       _ f p t o s t r             s i z e I n B y t e s   >   ( s i z e _ t ) ( ( d i g i t s   >   0   ?   d i g i t s   :   0 )   +   1 )                           p f l t   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ c o n v \ c f o u t . c                 _ f l t o u t 2         s t r c p y _ s ( r e s u l t s t r ,   r e s u l t s i z e ,   a u t o f o s . m a n )                         ( o p t i o n s   &   ~ _ T W O _ D I G I T _ E X P O N E N T )   = =   0                       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ o u t p u t f o r m a t . c                       _ s e t _ o u t p u t _ f o r m a t             ( " I n v a l i d   i n p u t   v a l u e " ,   0 )             f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ t r a n \ c o n t r l f p . c                   _ c o n t r o l f p _ s         �E N U   (�E N U   P�E N U   x�E N A   ��N L B   ��E N C   ��Z H H   ��Z H I   ��C H S   ��Z H H   �C H S   D�Z H I   p�C H T   ��N L B   ��E N U   ��E N A   �E N L   ,�E N C   H�E N B   t�E N I   ��E N J   ��E N Z   ��E N S   �E N T   H�E N G   d�E N U   ��E N U   ��F R B   ��F R C   ��F R L   �F R S   4�D E A   \�D E C   ��D E L   ��D E S   ��E N I   ��I T S    �N O R   8�N O R   `�N O N   ��P T B   ��E S S   ��E S B   �E S L   8�E S O   `�E S C   ��E S D   ��E S F   ��E S E   (�E S G   T�E S H   |�E S M   ��E S N   ��E S I   ��E S A   �E S Z   @�E S R   `�E S U   ��E S Y   ��E S V   ��S V F   �D E S   �E N G   �E N U   $�E N U                                                                                                                                                               a m e r i c a n         a m e r i c a n   e n g l i s h         a m e r i c a n - e n g l i s h         a u s t r a l i a n         b e l g i a n       c a n a d i a n         c h h       c h i       c h i n e s e       c h i n e s e - h o n g k o n g         c h i n e s e - s i m p l i f i e d             c h i n e s e - s i n g a p o r e           c h i n e s e - t r a d i t i o n a l           d u t c h - b e l g i a n           e n g l i s h - a m e r i c a n         e n g l i s h - a u s       e n g l i s h - b e l i z e         e n g l i s h - c a n       e n g l i s h - c a r i b b e a n           e n g l i s h - i r e       e n g l i s h - j a m a i c a           e n g l i s h - n z         e n g l i s h - s o u t h   a f r i c a             e n g l i s h - t r i n i d a d   y   t o b a g o               e n g l i s h - u k         e n g l i s h - u s         e n g l i s h - u s a       f r e n c h - b e l g i a n         f r e n c h - c a n a d i a n           f r e n c h - l u x e m b o u r g           f r e n c h - s w i s s         g e r m a n - a u s t r i a n           g e r m a n - l i c h t e n s t e i n           g e r m a n - l u x e m b o u r g           g e r m a n - s w i s s         i r i s h - e n g l i s h           i t a l i a n - s w i s s           n o r w e g i a n       n o r w e g i a n - b o k m a l         n o r w e g i a n - n y n o r s k           p o r t u g u e s e - b r a z i l i a n             s p a n i s h - a r g e n t i n a           s p a n i s h - b o l i v i a           s p a n i s h - c h i l e           s p a n i s h - c o l o m b i a         s p a n i s h - c o s t a   r i c a             s p a n i s h - d o m i n i c a n   r e p u b l i c             s p a n i s h - e c u a d o r           s p a n i s h - e l   s a l v a d o r           s p a n i s h - g u a t e m a l a           s p a n i s h - h o n d u r a s         s p a n i s h - m e x i c a n           s p a n i s h - m o d e r n         s p a n i s h - n i c a r a g u a           s p a n i s h - p a n a m a         s p a n i s h - p a r a g u a y         s p a n i s h - p e r u         s p a n i s h - p u e r t o   r i c o           s p a n i s h - u r u g u a y           s p a n i s h - v e n e z u e l a           s w e d i s h - f i n l a n d           s w i s s       u s     u s a       |�U S A   ��G B R   ��C H N   ��C Z E   ��G B R   ��G B R   ��N L D   �H K G   (�N Z L   D�N Z L   L�C H N   d�C H N   |�P R I   ��S V K   ��Z A F   ��K O R   ��Z A F   �K O R    �T T O   �G B R   L�G B R   p�U S A   �U S A                                                           a m e r i c a       b r i t a i n       c h i n a       c z e c h       e n g l a n d       g r e a t   b r i t a i n           h o l l a n d       h o n g - k o n g       n e w - z e a l a n d       n z     p r   c h i n a         p r - c h i n a         p u e r t o - r i c o       s l o v a k     s o u t h   a f r i c a         s o u t h   k o r e a       s o u t h - a f r i c a         s o u t h - k o r e a       t r i n i d a d   &   t o b a g o           u n i t e d - k i n g d o m         u n i t e d - s t a t e s           A          f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ g e t q l o c . c                   _ _ g e t _ q u a l i f i e d _ l o c a l e             w c s n c p y _ s ( l p O u t S t r - > s z L o c a l e N a m e ,   ( s i z e o f ( l p O u t S t r - > s z L o c a l e N a m e )   /   s i z e o f ( l p O u t S t r - > s z L o c a l e N a m e [ 0 ] ) ) ,   _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   w c s l e n ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   +   1 )                                                                           L a n g C o u n t r y E n u m P r o c E x           w c s n c p y _ s ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   ( s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   /   s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e [ 0 ] ) ) ,   l p L o c a l e S t r i n g ,   w c s l e n ( l p L o c a l e S t r i n g )   +   1 )                                                                         L a n g u a g e E n u m P r o c E x             G e t L o c a l e N a m e F r o m D e f a u l t             w c s n c p y _ s ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   ( s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   /   s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e [ 0 ] ) ) ,   l o c a l e N a m e ,   w c s l e n ( l o c a l e N a m e )   +   1 )                                                                     A C P       O C P       6-    ( p a t h   ! =   N U L L )             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ o p e n . c                   _ o p e n       ( p f h   ! =   N U L L )           _ s o p e n _ h e l p e r               ( ( p m o d e   &   ( ~ ( _ S _ I R E A D   |   _ S _ I W R I T E ) ) )   = =   0 )                     s 1   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m b s t r i n g \ m b s n b c m p . c                     _ m b s n b c m p _ l       s 2   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m b s t r i n g \ m b s n b i c m . c                     _ m b s n b i c m p _ l         _ w o p e n     _ w s o p e n _ h e l p e r         CreateFile2     _ w s o p e n _ n o l o c k         _ g e t _ f m o d e ( & f m o d e )             (   " I n v a l i d   o p e n   f l a g "   ,   0   )               (   " I n v a l i d   s h a r i n g   f l a g "   ,   0   )                     ( o f l a g   &   ( _ O _ T E X T   |   _ O _ W T E X T   |   _ O _ U 1 6 T E X T   |   _ O _ U 8 T E X T )   )   ! =   0                           0   & &   " I n t e r n a l   E r r o r "           0   & &   " O n l y   U T F - 1 6   l i t t l e   e n d i a n   &   U T F - 8   i s   s u p p o r t e d   f o r   r e a d s "                               f i r s t   ! =   N U L L           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ w c s n i c m p . c                     _ w c s n i c m p _ l       l a s t   ! =   N U L L         _ w c s n i c m p       _ o u t p u t _ p _ l       ( ( t y p e _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                 ( " I n c o r r e c t   f o r m a t   s p e c i f i e r " ,   0 )                       ( ( w i d t h _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                       _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ w i d t h _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                   ( ( p r e c i s _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                     _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ p r e c i s _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                 ( ( t y p e _ p o s > = 0 )   & &   ( t y p e _ p o s < _ A R G M A X ) )                       _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ s h o r t _ a r g ,   c h ,   f l a g s )                                 _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ p t r _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ d o u b l e _ a r g ,   c h ,   f l a g s )                               p a s s   = =   F O R M A T _ O U T P U T _ P A S S             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t 6 4 _ a r g ,   c h ,   f l a g s )                                 _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ l o n g _ l o n g _ a r g ,   c h ,   f l a g s )                                 ( ( s t a t e   = =   S T _ N O R M A L )   | |   ( s t a t e   = =   S T _ T Y P E ) )                         ( " M i s s i n g   p o s i t i o n   i n   t h e   f o r m a t   s t r i n g " ,   0 )                         ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp                       _ o u t p u t _ s _ l       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ p r i n t f . c                   p r i n t f     s i z e I n B y t e s   < =   I N T _ M A X             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ w c t o m b . c                   _ w c t o m b _ s _ l       ( o p t i o n   ! =   N U L L )         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ g e t e n v . c                     g e t e n v     ( _ t c s n l e n ( o p t i o n ,   _ M A X _ E N V )   <   _ M A X _ E N V )                   _ t c s n l e n ( * s e a r c h   +   l e n g t h   +   1 ,   _ M A X _ E N V )   <   _ M A X _ E N V                       p R e t u r n V a l u e   ! =   N U L L             _ g e t e n v _ s _ h e l p e r         ( b u f f e r   ! =   N U L L   & &   s i z e I n T C h a r s   >   0 )   | |   ( b u f f e r   = =   N U L L   & &   s i z e I n T C h a r s   = =   0 )                                       s t r c p y _ s ( b u f f e r ,   s i z e I n T C h a r s ,   s t r )                   p B u f f e r   ! =   N U L L           _ d u p e n v _ s _ h e l p e r         v a r n a m e   ! =   N U L L           s t r c p y _ s ( * p B u f f e r ,   s i z e ,   s t r )               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ t m a k e p a t h _ s . i n l                     _ w m a k e p a t h _ s         ( ( ( _ P a t h ) ) )   ! =   N U L L           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ t s p l i t p a t h _ s . i n l                       _ w s p l i t p a t h _ s           ( L " I n v a l i d   p a r a m e t e r " ,   0 )               C O N O U T $       _ w o u t p u t _ p _ l         _ w o u t p u t _ s _ l             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f p u t w c . c                   f p u t w c     _ L o c a l e   ! =   N U L L           f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ i n c l u d e \ s t r g t o l d 1 2 . i n l                     _ _ s t r g t o l d 1 2 _ l             f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ c o n v \ x 1 0 f o u t . c                     $ I 1 0 _ O U T P U T           s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # S N A N " )                 1#SNAN      s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N D " )                   1#IND       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N F " )                   1#INF       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # Q N A N " )                 1#QNAN   f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ t r a n \ i 3 8 6 \ i e e e 8 7 . c                     _ s e t _ c o n t r o l f p             _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   n e w c t r l ,   m a s k   &   ~ 0 x 0 0 0 8 0 0 0 0 )                             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ s t r n i c m p . c                     _ s t r n i c m p _ l       c o u n t   < =   I N T _ M A X         _ s t r n i c m p           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ c h s i z e . c                   _ c h s i z e _ s       ( s i z e   > =   0 )           ( ( m o d e   = =   _ O _ T E X T )   | |   ( m o d e   = =   _ O _ B I N A R Y )   | |   ( m o d e   = =   _ O _ W T E X T )   | |   ( m o d e   = =   _ O _ U 8 T E X T )   | |   ( m o d e   = =   _ O _ U 1 6 T E X T ) )                                                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ s e t m o d e . c                     _ s e t m o d e             ( ( m o d e   = =   _ O _ T E X T )   | |   ( m o d e   = =   _ O _ B I N A R Y )   | |   ( m o d e   = =   _ O _ W T E X T ) )                             _ s e t _ f m o d e         ( p M o d e   ! =   N U L L )           _ g e t _ f m o d e         n p t r   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ s t r t o l . c                   s t r t o x l       i b a s e   = =   0   | |   ( 2   < =   i b a s e   & &   i b a s e   < =   3 6 )                       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ v p r i n t f . c                     v p r i n t f _ h e l p e r         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ s t r t o q . c                   s t r t o x q       f:\dd\vctools\crt\crtw32\misc\wtombenv.c                f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m b s t r i n g \ m b s n b i c o . c                     _ m b s n b i c o l l _ l           n   < =   I N T _ M A X         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ w c s t o l . c                   w c s t o x l       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ w c s t o q . c                   w c s t o x q       f:\dd\vctools\crt\crtw32\convert\wcstoq.c               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ s t r t o d . c                   _ s t r t o d _ l       p o p t i o n   ! =   N U L L               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ s e t e n v . c                     _ _ c r t s e t e n v       e q u a l   -   o p t i o n   <   _ M A X _ E N V                   _ t c s n l e n ( e q u a l   +   1 ,   _ M A X _ E N V )   <   _ M A X _ E N V                     f:\dd\vctools\crt\crtw32\misc\setenv.c              ( " C R T   L o g i c   e r r o r   d u r i n g   s e t e n v " , 0 )                   s t r c p y _ s ( n a m e ,   s t r l e n ( o p t i o n )   +   2 ,   o p t i o n )                     c o p y _ e n v i r o n         s t r c p y _ s ( * n e w e n v p t r ,   e n v p t r S i z e ,   * o l d e n v p t r )                     _ s t r i n g 1   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ s t r n i c o l . c                     _ s t r n i c o l l _ l         _ s t r i n g 2   ! =   N U L L         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ w c s t o d . c                   _ w c s t o d _ l       s t r i n g   ! =   N U L L         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m b s t r i n g \ m b s c h r . c                     _ m b s c h r _ l       _ _ w s t r g t o l d 1 2 _ l           H                                                           ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                RSDS�)?��E�N�ww�4d   C:\Program Files\MAXON\CINEMA 4D R13\plugins\STL_Importer\obj\STL_Importer_Win32_Debug.pdb      ;  ;                                                                                                                                                                                                                                                                                                     H�        ����    @   P                   d    ,                ��               �    ��    �       ����    @   �        (�        ����    @   �                         �                D�                 4     @ d     D�       ����    @             d�       ����    @   �                    �     �     d�        ����    @   �                     ���                �     !@ d     ��       ����    @   �                     ��@!               T!    \!    ��        ����    @   @!                  ��!               �!    �!�!","    �       ����    @   �!        ��              P   �         D�              @             d�              @   �                     X�h"               |"    �"\!    X�       ����    @   h"            p      ���"               �"    �"�!�!","        ��       ����    @   �"                     �0#               D#    P#,     �       ����    @   0#                    ���#               �#    �#    ��        ����    @   �#        �       ����    @   �#                   $    �#�#                ��#                4�@$               T$    d$�#�#    4�       ����    @   @$                    \��$               �$    �$�#�#    \�       ����    @   �$                    �� %               %    (%�$�#�#    ��       ����    @    %                    ��d%               x%    �%    ��        ����    @   d%                    ���%               �%    �%P#,    ��       ����    @   �%                    ��&               0&    D&�%P#,    ��       ����    @   &                    ���&               �&    �&�%    ��       ����    @   �&                     ��&               �&     '�&�%     �       ����    @   �&                    4�<'               P'    `'�&�%    4�       ����    @   <'                    l��'               �'    �'D&�%P#,        l�       ����    @   �'                    h�(               (    0(d$�#�#    h�       ����    @   (                    ��l(               �(    �(��    ��       ����    @   l(                    (��                ���(               �(     )    ��        ����    @   �(                    ��<)               P)    X)    ��        ����    @   <)                    ���)               �)    �)X)    ��       ����    @   �)                    ��)               *    *    �        ����    @   �)                    8�H*               \*    d*    8�        ����    @   H*                    X��*               �*    �*    X�        ����    @   �*                    |��*               +    +X)    |�       ����    @   �*                    ��T+               h+    t+,    ��       ����    @   T+                    ���+               �+    �+,    ��       ����    @   �+                    ��,                ,    0,�+,    ��       ����    @   ,                    �l,               �,    �,�+,    �       ����    @   l,                    @��,               �,    �,�+,    @�       ����    @   �,                    h�,-               @-    P-P#,    h�       ����    @   ,-                    ���-               �-    �-,    ��       ����    @   �-                    ���-               �-    .P#,    ��       ����    @   �-                    ��H.               \.    l.�#�#    ��       ����    @   H.                    ��.               �.    �.�#�#    �       ����    @   �.                    p�/               /    ,/�#�#    p�       ����    @   /                    ��h/               |/    �/�#�#    ��       ����    @   h/                    ���/               �/    �/d$�#�#    ��       ����    @   �/                    $�,0               @0    T0d$�#�#    $�       ����    @   ,0                    L��0               �0    �0�$�#�#    L�       ����    @   �0                    p��0               1    1�$�#�#    p�       ����    @   �0                    ��X1               l1    |1�#�#    ��       ����    @   X1                     ��1               �1    �1�#�#     �       ����    @   �1                    d�2               ,2    <2�#�#    d�       ����    @   2                    ��x2               �2    �2�#�#    ��       ����    @   x2                    ���2               �2    �2�#�#    ��       ����    @   �2                    ��83               L3    \3�#�#    ��       ����    @   83                     ��3               �3    �3�#�#     �       ����    @   �3                    h��3               4    4�#�#    h�       ����    @   �3                    ��X4               l4    �4�2�#�#    ��       ����    @   X4                    ���4               �4    �4�#�#    ��       ����    @   �4                     �5               05    @5�#�#     �       ����    @   5                    ��|5               �5    �5�5�2�#�#        ��       ����    @   |5        ��       ����    @   �5                   6    �5�2�#�#                ��46               H6    d6�5�2�#�#        ��       ����    @   46                    ��6               �6    �6\3�#�#    �       ����    @   �6                    x�7               7    (7�#�#    x�       ����    @   7                    ���5                ��|7               �7    �7�#�#    ��       ����    @   |7                    D��7               �7     8�#�#    D�       ����    @   �7                    l�<8               P8    `8�#�#    l�       ����    @   <8                    ���8               �8    �8�2�#�#    ��       ����    @   �8                    �� 9               9    $9�#�#    ��       ����    @    9                     �`9               t9    �9�#�#     �       ����    @   `9                    ���9               �9    �9:�2�#�#        ��       ����    @   �9        ��       ����    @   8:                   L:    :�2�#�#                ��x:               �:    �::�2�#�#        ��       ����    @   x:                     ��:               �:    ;\3�#�#     �       ����    @   �:                    h�H;               \;    l;�#�#    h�       ����    @   H;                    ��8:                ���;               �;    �;�#�#    ��       ����    @   �;                    �� <               4<    H<�2�#�#    ��       ����    @    <                    ��<               �<    �<�#�#    �       ����    @   �<                    ���<               �<    =�#�#    ��       ����    @   �<                    ��D=               X=    t=�=�2�#�#        ��       ����    @   D=        �       ����    @   �=                   �=    �=�2�#�#                4��=               >    ,>�=�2�#�#        4�       ����    @   �=                    `�h>               |>    �>\3�#�#    `�       ����    @   h>                    ���>               �>    �>�#�#    ��       ����    @   �>                    ��=                H�P                ��\?               p?    |?,    ��       ����    @   \?                    ,��?               �?    �?,    ,�       ����    @   �?                    P�@               (@    8@�?,    P�       ����    @   @                    |�t@               �@    �@    |�        ����    @   t@                    ���@               �@    �@,    ��       ����    @   �@                    ��(A               <A    DA    ��        ����    @   (A                    ���A               �A    �ADA    ��       ����    @   �A                    ���A               �A    �ADA    ��       ����    @   �A                    �8B               LB    XBDA    �       ����    @   8B                    4��B               �B    �BDA    4�       ����    @   �B                    X��B               C    CDA    X�       ����    @   �B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �{	            |	����    ����                  "�   @L   �L                            0L               L                            ��	����    ����                  �L"�   �L   �L                                    ��	����    ����                  M"�   ,M   <M                                    #�	����    ����                  |M"�   �M   �M                                    *	����    ����                  �M"�   �M   �M                                    �	����    ����                  <N"�   LN   \N                                    �����    ����                  �N"�   �N   �N                                    �����    ����                  �N"�   O   O                            �(    pO       �O�O         �    ����       MF        H�    ����       i        �Q    �O       �OP0P�O�O        l�    ����       7        ��    ����       �I        ��    ����       =        U*    dP       tP�O        ��    ����       <C        Q$    �P       �P�O       ��    ����       r]        �n    �P        Q Q�O        ��    ����       L        ��    ����       P        6&    TQ       hQ Q�O        �    ����       �C        �R    �Q       �Q Q�O        @�    ����       �E        ?    �Q       �Q�O�O        h�    ����       �D        wg    ,R       <R�O        ��    ����       �h        $`    pR       �R�O�O        ��    ����       �;    ���� �"�   �R                           �����"�   �R                           ������"�   S                           ������"�   4S                           ������"�   dS                           ������    ��"�   �S                               ����@�    H�"�   �S                               ����P�"�   T                           ������������"�   <T                               "�   �T                       ��������������������������� �        ���� �    �"�   �T                               ����0�    K�����K�"�   U                               ����0�"�   LU                           "�   �U                       ����@�����K�   S�   ^�����f�        ������"�   �U                           ������"�    V                           ���� �"�   0V                           ����@�"�   `V                           ������"�   �V                           ���� �"�   �V                           ������"�   �V                           ����`�    h�"�    W                               ������������   ��   ��"�   \W                               ������������   �   �"�   �W                               ������"�   �W                           ������    ��������"�   $X                               ����`�"�   hX                           ������������"�   �X                               ������������   ��   ��"�   �X                               ������������    �   �"�    Y                               ������"�   lY                           ������"�   �Y                           �����    +�����+�"�   �Y                               @           Dy����    ����                  Z"�    Z   0Z                       ���� �"�   pZ                           ����`�"�   �Z                           "�   �Z                       ��������������������������������������������:�����U�����p�������������������                "�   �[                       ����������������������������	�����$�����?�����Z�����u�������������������������                ����@"�   \                           ������"�   8\                           ������    ��������"�   h\                               ������"�   �\                           ���� �    ;�����;�"�   �\                               ����p�"�    ]                           ������    ��������"�   P]                               ����@�"�   �]                           ���� �    ;�����;�"�   �]                               ������"�   ^                           ����`�"�   8^                           �����"�   h^                           ������"�   �^                           ����P�"�   �^                           ���� �"�   �^                           ������"�   (_                           ������"�   X_                           "�
   �_                       ����0    8   @   H   P   X   c   k   v   �            @           �K@           %L����    ����                  "�   (`   l`                           `              `                ������    ��"�   �`                               ������    ��"�   �`                               ����0�    K�����K�"�   a                               ������"�   `a                           ����P    X"�   �a                               ������    ��������"�   �a                               ������"�   b                           "�   db                       ����0 ����;    C    N ����V         ����p�"�   �b                           ������"�   �b                           ������"�   �b                           ����0�"�   $c                           ������"�   Tc                           ������"�   �c                           ����p�"�   �c                           �����    �"�   �c                               ����������   #�   .�"�    d                               ������������   �   �"�   ld                               ������"�   �d                           ������    ��������"�   �d                               ����P�"�   ,e                           ����������"�   \e                               ������������   ��   ��"�   �e                               ����@�����H�   P�   X�"�   �e                               ����0�"�   0f                           ������"�   `f                           ����p�    ��������"�   �f                               @           �����    ����                  �f"�   �f   �f                       ������"�   4g                           �����"�   dg                           "�   �g                       ������    ��   ��������   ��        �����    �    "�   �g                               ����0�"�   ,h                           ������"�   \h                           ����`�    x�����x�"�   �h                               ������"�   �h                           ����0�"�    i                           ����0�    K�����K�"�   0i                               ������"�   ti                           ���� �"�   �i                           "�   �i                       ����P�����[�����f�   n�   v�   ��   ��   ��   ��   ��   ��
   ��   �   2�   T�   _�   g�   r�   }�   ��                    ����P�"�   �j                           ������"�   �j                           �����    +�����+�"�   k                               ��������"�   Pk                               ����������"�   �k                               "�   �k                       ����@�    H�    S�    ^�   f�   n�   v�   ��   ��   ��   ��   ��   ��   ��   ��                �����"�   tl                           ������"�   �l                           ������"�   �l                           @           ������    ����                  m"�   m   $m                       ������    ��������"�   dm                               ����p�"�   �m                           ����`�    {�����{�"�   �m                               ����@�"�   n                           �����"�   Ln                           ����P�    k�����k�"�   |n                               @           8����    ����                  �n"�   �n   �n                       �����"�    o                           ����0"�   Po                           �����"�   �o                           ����� "�   �o                           ������"�   �o                           ������"�   p                           ����P�"�   @p                           ������"�   pp                           ����@�    [�����[�"�   �p                               ������"�   �p                           "�   8q                       ���� ������   �   �����&�        ����@�"�   hq                           ������"�   �q                           ������"�   �q                           ���� �"�   �q                           ������"�   (r                           ������"�   Xr                           ����@�"�   �r                           ������    ��"�   �r                               ������������   ��   ��"�   �r                               ������������   ��   ��"�   @s                               ������"�   �s                           ���� �    ;�����;�"�   �s                               ���� �"�    t                           ����`����k"�   0t                               ����@�����K�   S�   ^�"�   lt                               ������������   ��   ��"�   �t                               ���� �"�   u                           ������"�   4u                           ���� �    ������"�   du                               @           �����    ����                  �u"�   �u   �u                       ����`�"�   v                           ������"�   8v                           "�   �v                       ���� �    �   1������   1�        �����    �   �"�   �v                               ���� �"�    w                           ������"�   0w                           ���� �    ������"�   `w                               ������"�   �w                           ���� �"�   �w                           ������    ��������"�   x                               ����@�"�   Hx                           ������"�   xx                           "�   �x                       ����`�����k�����v�   ~�   ��   ��   ��   ��   ��   ��   ��
   ��    �   B�   d�   o�   w�   ��   ��   ��                    ���� �"�   �y                           ����`�"�   �y                           ������    ��������"�   �y                               ����p����x"�   $z                               ���� ����("�   `z                               "�   �z                       ����@�    H�    S�    ^�   f�   n�   v�   ��   ��   ��   ��   ��   ��   ��   ��                ������"�   H{                           ������"�   x{                           ����`�"�   �{                           ����0�"�   �{                           ���� �"�   |                           ������"�   8|                           "�
   �|                       �����    �   �   �   �   �   �   �   �   �            @           �I@           �I����    ����                  "�   }   L}                           �|              �|                ����`�    h�"�   �}                               ������"�   �}                           ������"�   �}                           ������"�    ~                           @           ������    ����                  P~"�   `~   p~                       ������    ������"�   �~                               �����"�   �~                           ������    ��������"�   $                               ������"�   h                           ������"�   �                           ������    ��������"�   �                               @           X����    ����                  �"�   �   ,�                       ����`"�   l�                           ���� "�   ��                           �����"�   ̀                           ����� "�   ��                           ����`�"�   ,�                           ������"�   \�                           ����@�    H�"�   ��                               ������    ��������"�   ȁ                               ������"�   �                           ����     "�   <�                               ���� �"�   x�                           ������"�   ��                           ����p�"�   ؂                           ������"�   �                           ���� �"�   8�                           ����P�"�   h�                           ���� �"�   ��                           ������"�   ȃ                           ����@�"�   ��                           ������"�   (�                           ������"�   X�                           ������"�   ��                           ������"�   ��                           ����@�"�   �                           "�	   <�                       ������    ��   ��   ��   ��   ��   ��   ��   ��            "�	   ��                       ����@�    H�   P�   X�   `�   h�   p�   `�   p�            ����`�"�   �                           ���� �"�   8�                           �����"�   h�                           "�
   ��                       ����0    8   @   H   P   X   c   k   v   �            ����@    H"�   �                               "�   x�                       ���� ����8����P����h��������������������            ���� 	"�   ć                           "�   �                       �����
    �
   �����
           �����    �   �"�   H�                               ����@"�   ��                           ����P	"�   ��                           ����p    ������"�   �                               ����p"�   0�                           �����	"�   `�                           �����    ������"�   ��                               �����"�   ԉ                           �����"�   �                           "�   X�                       ���������������   �   �   �   �   �   �      
   >   `   �   �   �   �   �   �   �                    �����"�   �                           �����	"�   <�                           ����@    [����["�   l�                               ����@����H"�   ��                               ����������"�   �                               "�   L�                       �����    �    �    �   �   �   �   �   �            (   3   >                �����"�   Ԍ                           �����"�   �                           �����"�   4�                           @           �{����    ����                  d�"�   t�   ��                       ����     ;����;"�   č                               ����0"�   �                           �����    ������"�   8�                               ���� "�   |�                           �����	"�   ��                           �����    ������"�   ܎                               @           X~����    ����                   �"�   0�   @�                       �����"�   ��                           ����`"�   ��                           �����"�   ��                           ����0"�   �                           ����p"�   @�                           ����`"�   p�                           ����
    
"�   ��                               ����     ����"�   ܐ                               �����"�    �                           �����    �"�   P�                               �����"�   ��                           �����
"�   ��                           ����P
"�   �                           �����
"�   �                           "�	   p�                       �����    �   �   �   �   �       �                    ����    ����    ����    �a    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    R�        %�        ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    '�    ����    ����    ����    7�    ����    ����    ����    Π    ����    ����    ����    ��    ����    ����    ����    ?�    ����    ����    ����    ��    ����    ����    ����    =�    ����    ����    ����    '�    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    I�    ����    ����    ����    !�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    O�    ����    ����    ��������    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����*    ����    ����    ����    "    ����    ����    ����    [C    +C8C        ����    ����    ����    Y'    _&l&        ����    ����    �����6�6    ����    ����    �����#$    @           
)����    ����                  �"�   (�   8�                       ����    ����    ����	::        �5    ��       ���O        ��    ����       <H        ����    ����    ����    {g    ����    ����    ����    �j    ����    ����    ����    
o    ����    ����    ����    �r    ���� "�   `�                           ����    ����    ��������    ����    ����    ��������    ����    ����    ����    5    ����    ����    ����%4U4    ����    ����    ����    #A    ����    ����    ����    �E    ����    ����    ����    �H    ����    d���    ����    >b    ����    ����    ����    Ze    ����    ����    ����    �t    ����    ����    ����    fx    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    �        W�        ����    ���    ����    ��        ʤ        ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    a�    ����0"�   �                           ����    ����    ����    =�    ����    ����    ����    ������    �        ����    ����    ����    ������    3�        ����    ����    ����W�]�    ����    ����    ��������    ����    ����    ����    s�    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    q�    ����    ����    ����    r�    ����    ����    ����    �0����    �0        ����    ����    ����    �.����    Z/        ����    ����    ����    Z6        _5        '6            ����    ����    ����    �     ����    ����    ����    b    ����    ����    ����    �w    ����    ����    ����    Vz    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ��������    ����    ����    ����             �        ����    ����    ����        ����    ����    ����    �    ����    ����    ����        ����    ����    ����    }    ����    |���    ����    r    ����    |���    ����    (s    ����`"�   P�                           ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    5�    ����    ����    ����    ��    ����    ����    ����    �U    ����    ����    ����    �_    ����    ����    ����    4g    ����    ����    ����    1h    ����    ����    ����    :�    ����    ����    ����    �)    ����    ����    ����    /    �����"�   �                           ����    ����    ����    8<    �����"�   0�                           ���� "�   `�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               P�Z    ��          �� �� �� fP ��   STL_Importer.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �   8   �   �      ^  �  B  �  Q   �   �   �  �  �   D   g   �   -   ����       
       Copyright (c) 1992-2004 by P.J. Plauger, licensed by Dinkumware, Ltd. ALL RIGHTS RESERVED.                                       �              �             �               3              �9               A                                         �              �              �             �              �<              @>              2@                                             �              �             �              �<              @>              2@                                `�    `�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             t���������      ����        N�@���Du�  s�                  sqrt                                                                                                                                                                                                                                                                                                                                                         8�:�    ����   (�.   $�t�t�t�t�t�t�t�t�t�x�x�x�x�x�x�x�x�.                                                        	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                    zU          �      ���������              �           @]   D]   H]   L]   T]   \]!   d]   l]   t]   |]   �]   �]   �]   �]    �]   �]   �]   �]   �]   �]   �]   �]   �]   �]"   �]#   �]$   �]%   �]&   �]                                                       �D        � 0                �����
                                                                               ����������������                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                                     abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                            X��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                                                                                                                            P����   C   ܁���������� ��� �,�4�@�D�H�L�P�T�X�\�`�d�h�l�p�|�����P�����������ȂԂ������       �$�0�<�H�T�`�l�|�������Ѓ�������(�4�@�L�X�d�p�|�������Ą(�Ԅ������(�@�X�`�h�����`                                                                        8�                                   ��            ��            ��            ��            ��                          (�        8���@���                                                            8�X�    ����            �T�T�T�T�T�T�T�T�T�T        <�            ���    ����        ����            �p     ����    PST                                                             PDT                                                             ����                                �&                                                                                                                                                                                                                                                                       �                            ����   :   Y   w   �   �   �   �     /  M  l  ����   ;   Z   x   �   �   �   �     0  N  m                      ����   ���5      @   �  �   ����                                      �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                                          �                                                                                                                                                                                                                                                                                                                                                        ��    .?AVruntime_error@std@@         ��    .?AVexception@std@@         ��    .?AVfailure@ios_base@std@@          ��    .?AVsystem_error@std@@          ��    .?AV_System_error@std@@         ��    .?AVbad_cast@std@@      ��    .?AVCommandData@@       ��    .?AVBaseData@@      ��    .?AVios_base@std@@      ��    .?AV?$_Iosb@H@std@@         ��    .?AV?$basic_ios@DU?$char_traits@D@std@@@std@@           ��    .?AV?$basic_streambuf@DU?$char_traits@D@std@@@std@@             ��    .?AV?$basic_istream@DU?$char_traits@D@std@@@std@@               ��    .?AV?$basic_filebuf@DU?$char_traits@D@std@@@std@@               ��    .?AV?$basic_ifstream@DU?$char_traits@D@std@@@std@@              ��    .?AV_Facet_base@std@@       ��    .?AVfacet@locale@std@@          ��    .?AVcodecvt_base@std@@          ��    .?AUctype_base@std@@        ��    .?AV?$ctype@D@std@@         ��    .?AVerror_category@std@@        ��    .?AV_Generic_error_category@std@@           ��    .?AV_Iostream_error_category@std@@          ��    .?AV_System_error_category@std@@            ��    .?AV?$codecvt@DDH@std@@         ��    .?AVSimplePlugin@@      ��    .?AVNeighbor@@      ��    .?AVGeSortAndSearch@@       ��    .?AVDisjointNgonMesh@@          ��    .?AVGeToolNode2D@@      ��    .?AVGeToolList2D@@      ��    .?AVGeToolDynArray@@        ��    .?AVGeToolDynArraySort@@        ��    .?AVbad_alloc@std@@         ��    .?AVinvalid_argument@std@@          ��    .?AVlogic_error@std@@       ��    .?AVlength_error@std@@          ��    .?AVout_of_range@std@@          ��    .?AVoverflow_error@std@@        ��    .?AVbad_function_call@std@@         ��    .?AVregex_error@std@@       ��    .?AV_Locimp@locale@std@@        ��    .?AV?$num_get@DV?$istreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                       ��    .?AV?$num_put@DV?$ostreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                   ��    .?AV?$numpunct@D@std@@          ��    .?AV?$codecvt@_WDH@std@@        ��    .?AV?$codecvt@GDH@std@@         ��    .?AV?$ctype@_W@std@@        ��    .?AV?$ctype@G@std@@             ��    .?AV?$num_get@_WV?$istreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                    ��    .?AV?$num_get@GV?$istreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                   ��    .?AV?$numpunct@_W@std@@         ��    .?AUmessages_base@std@@         ��    .?AUmoney_base@std@@        ��    .?AUtime_base@std@@             ��    .?AV?$num_put@_WV?$ostreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                    ��    .?AV?$collate@_W@std@@          ��    .?AV?$messages@_W@std@@         ��    .?AV?$money_get@_WV?$istreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                  ��    .?AV?$money_put@_WV?$ostreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                  ��    .?AV?$moneypunct@_W$0A@@std@@           ��    .?AV?$_Mpunct@_W@std@@          ��    .?AV?$moneypunct@_W$00@std@@            ��    .?AV?$time_get@_WV?$istreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                   ��    .?AV?$time_put@_WV?$ostreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                   ��    .?AV?$num_put@GV?$ostreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                   ��    .?AV?$numpunct@G@std@@          ��    .?AV?$collate@G@std@@       ��    .?AV?$messages@G@std@@          ��    .?AV?$money_get@GV?$istreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                     ��    .?AV?$money_put@GV?$ostreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                 ��    .?AV?$moneypunct@G$0A@@std@@        ��    .?AV?$_Mpunct@G@std@@       ��    .?AV?$moneypunct@G$00@std@@         ��    .?AV?$time_get@GV?$istreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                      ��    .?AV?$time_put@GV?$ostreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                  ��    .?AV?$collate@D@std@@       ��    .?AV?$messages@D@std@@          ��    .?AV?$money_get@DV?$istreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                     ��    .?AV?$money_put@DV?$ostreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                 ��    .?AV?$moneypunct@D$0A@@std@@        ��    .?AV?$_Mpunct@D@std@@       ��    .?AV?$moneypunct@D$00@std@@         ��    .?AV?$time_get@DV?$istreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                      ��    .?AV?$time_put@DV?$ostreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                  ��    .?AVbad_typeid@std@@        ��    .?AV__non_rtti_object@std@@         ��    .?AVtype_info@@     ��    .?AVbad_exception@std@@         ��    .?AVDNameNode@@     ��    .?AVcharNode@@      ��    .?AVpcharNode@@     ��    .?AVpDNameNode@@        ��    .?AVDNameStatusNode@@       ��    .?AVpairNode@@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  � � �    0 F \ n � � � � � � �   0 @ L h � � � � � � � 
  & 0 B R f x � � � � � � �   0 B R ^ l ~ � � � � � � �   6 F \ l ~ � � � � � � � �   4 J d ~ � � � � � � �                                                                                                                  �         (                       � � �    0 F \ n � � � � � � �   0 @ L h � � � � � � � 
  & 0 B R f x � � � � � � �   0 B R ^ l ~ � � � � � � �   6 F \ l ~ � � � � � � � �   4 J d ~ � � � � � � �                                                                                                                  %EnterCriticalSection  �LeaveCriticalSection  DeleteCriticalSection !EncodePointer � DecodePointer �WideCharToMultiByte �MultiByteToWideChar �GetStringTypeW  gIsDebuggerPresent mIsProcessorFeaturePresent cGetModuleFileNameW  fGetModuleHandleExW  ;HeapValidate  �GetSystemInfo @RaiseException  �RtlUnwind �GetCommandLineA GetCurrentThreadId  XFatalAppExitA �GetCPInfo �UnhandledExceptionFilter  CSetUnhandledExceptionFilter SetLastError  HInitializeCriticalSectionAndSpinCount � CreateEventW  RSleep 	GetCurrentProcess aTerminateProcess  sTlsAlloc  uTlsGetValue vTlsSetValue tTlsFree �GetStartupInfoW �GetTickCount  gGetModuleHandleW  �GetProcAddress  � CreateSemaphoreW  PGetLastError  GetDateFormatW  �GetTimeFormatW  � CompareStringW  �LCMapStringW  TGetLocaleInfoW  tIsValidLocale �GetUserDefaultLCID  GEnumSystemLocalesW  �LoadLibraryExW  �GetStdHandle  �WriteFile QExitProcess  AreFileApisANSI  CloseHandle �FlushFileBuffers  �GetConsoleCP  �GetConsoleMode  >GetFileType PReadFile  �SetFilePointerEx  �SetConsoleCtrlHandler �OutputDebugStringW  �WaitForSingleObjectEx � CreateThread  �OutputDebugStringA  �WriteConsoleW rIsValidCodePage �GetACP  �GetOEMCP  3HeapFree  6HeapReAlloc 8HeapSize  5HeapQueryInformation  bGetModuleFileNameA  GetCurrentThread  /HeapAlloc �GetProcessHeap  -QueryPerformanceCounter 
GetCurrentProcessId �GetSystemTimeAsFileTime 'GetEnvironmentStringsW  �FreeEnvironmentStringsW �GetTimeZoneInformation  �VirtualQuery  �FreeLibrary "SetStdHandle  NReadConsoleW  � CreateFileW �SetEndOfFile  �SetEnvironmentVariableA KERNEL32.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                                             � (   �;	<_<i<�<�<!=q=�=>a>1?;?E?�?�? �   040>0d0n0�0�0�0�0�0161V1�1�1�1�1�1$2.2V2v2�2�2�2�2363V3t3�3�34444>4d4n4�4�4�4�455d5n5�5�5�5�5$6.6T6^6�6�6�6�6�6$7.7T7^7�7�7�7�7�78T8^8�8�8�8�8�89&9F9f9�9�9�9�9:&:F:f:�:�:�:�:;&;F;f;�;�;�;�;$<.<T<^<�<�<�<�<�<=6=V=v=�=�=�=�=>T>^>�>�>�>�>�>?&?F? � H   S0�4�4]5�5O6�6�7_;x;�;�;�;<_<x<�<�<�<�<G=`=l=�=W>�>�>?7?h?t?   �    v1�1�1�1I2v3�3�3�3I4  	 <   o0�0�0�0�0�0G1t1�1�12#2+2r2�2�2�23 3,30=�=�=�>8?\? 	 0   00�1�3D4v5�5<6`708�8�8;9H:�: ;v<�<?�?  	 $   0t0�0H1@2�2>3�3�5%6�6d9�9�? 0	 4   C0�0C1�1x2�2K45�56<6H6�9�9X:�:H;�>(?X?d?   @	 T   e2o2t2�2�3�3�3�3�344�5�5�5�5�5�5�5�5�5777 7%7.7G7L7Q7N8S8`8m8r8{8�8�8�8 P	 @   525y5 6�6�:�:�:+;5;�;�;<$<0<<<H<T<`<l<x<�<�<�<�<�<"?   `	 @   �023�3�4�4�45D5Y5|5�5�7�7�7�7�7818H8�;=�=�=�=�=?   p	 \   ~0�0Y1p1�2�2{314�4�4�4�4q5�5�5�5a6�6�6�6;:@:M:Z:_:k:�:�:�:�: ;<-<�<�<�<>3>d>p>�>   �	 (   M1|1�1�13J3x3�3�3*4X4d4�4647�? �	 8   �2505�6�647@7�8�:�:;$;�;�;a<�<= =v=�=$>�?�?   �	    >0$8�8�8�>? �	 $   0�0o1�1�3i4�4�8<,<b<r<�<�< �	    �4�4�6�7�89�?   �	     30`0l0?1�4�9:�:D<�<�<? �	 @   �2�2�2�2�2�24�4�4�4�5A6k6h8�8�8�8�8�8�8�8�8�899�?�?�? �	 0   �01H1T1�2M3T3�3�3�3d4k4�4k5r5�5�5�5�6�6  
 0   �0�1�4�4�4�4�4�4 57�7�7�7�:�;0<<<�?�?   
 T   �1�1�23�3�3�4"5�5s6�6�6�6�7�7U8�8�9�9�9�9�:�:e;<<<H<T<==�=�=�=>�>+?�?    
 \   0�01"1+1�13�3�3@4�4�56$606<6�6�7 8,888D89^:�:�:�:�:_;�;�;�<�<@=u= >?>�><?m?�?   0
 d   V0�001a1�1!2�2�233�3�3�3=4B4�45�5�5f6&7�7
8o8<9�9 :�:�:�:R;�;�;�;<?<�<K=�=V>�>�>?u?�?�? @
 X   �0�1�1�1�263\3�3�34<4�4�455"5/5�5�5�6
7=8�89�9:�:�:T;�;6<�<#=E=�=�=�>�>3?�? P
 T   /0�0/1�1V2�2�2�23�3�3U4�455�5o6�6[7�748�89�9=:�:';�;<�<=�=>�>�>v?�?   `
 H   V0�1�1�1:2�2"3�3
4z4�4]5�5]6�6�6�7i8]9�9;:�:2;�;4<�<"=?>�>.?�?   p
 P   D0�0$1�12t2�2�324�45�5�5d6�6�78�8K9p9|9�9R:�:�;�;k<�<O=�=�>�>�>;?�?   �
 L   60�01�1�2;3�34�4�56�6�6o7�7+9�9:+;�;�;�;<�<�<�<K=�=+>�>?{?�?   �
 L   [0�0;1�12�23�3�3{4�4_5�5R6�6K7�7?8�8$9�9:�:�:w;k<�<i=�=\>�>??�?   �
 D   �0/1�172�2/3{4�4s5�5K7�7+8�89�9�:Q;�;=�=�=�=C>h>t>�>k?�?   �
 L   L0�0+1�12{2�2\3�37'717;7E7O7Y7c7m7w7�7�7�7�7�7�7�7�;�;�;z=�=R>�>   �
 H   �1�2R3�3/4�4�4g5�5G6�6;7�7+8�8+9�9:x:�:x;�<�<�<K=�=>�>�>o?�?   �
 P   o0�0]1�1E2�2[3t4�4�4%5�5�677/8T8`8�8?9�9:�:�:k;�<�<�<+=�=>�>|?�?�?�? �
 L   k0�0K1o2�2�2�3�3 4/5T5`5�6�6�6�788�8�8k9�9[:t;�;�;<�<=/>T>`>�>W? �
 H   0^2�2K3�3B4�4G5�5;6�6+7[7�8�8�8�8�9�9::�:�;<�<�<V=�=N?�?�?     @   0 0,0�0{12�2�2�2�2�2m3�3a4�4a5�57�78�89�9�:O;J=>�>  8   �4O5�6�6_7�7T869�97:�:�:_;�;b<�<g=;>`>l>�>F?�?     `   /0�01�1�1t23�34v4�4]5�5/6�687�788�8:9�9:�:�:�:�:;�;�;�;<D<J<p<�<�<==�=?>�>9?�?   0 T   B0�0�01 1v1�1Y2�2�34o4�4V5�5M6�6&7�7)8�89}9�9?:�:;�;�;f<�<[=�=J>�>&?�?   @ h   
0z0�0V1�1B2�2"344�4�5�5�5V687\7h7�7W8�8�8�8�8�869�9�9::�:;;�;�;�;�;�;�;k<�<f=�=k>�>]?�?   P \   F0�0�01 1,181�12�23�3>4t4�4�4�4f5�5m6?7d7p7?8d8p8�8J9�9R:�:M;�;+<�<=�=�=}>�>e?   ` P   00�0Z1�1F2�2&3�34v4�4]5�5�6O7�7O8�89�9�9i:;�;<}<= =�>?Z?i?y?�?   p @   �0�01r2�2f3�3�4/5�5O6�6,7�768�8*9�9n:�:o;�<�< ==�?�?�? � X   60;0J0�0�0�0444!4.434S56666!6&6�9�9:L:Q:g:�;�;�<�<�=$>0><>H>T>`>�>�>�>�> � 4   z3�3h4�4f5�5V6�6c7�7m8�8[9K<�<?=�=/>�>[?�?   � D   {0�0m1�1b2�2]3�3;4�4>5�6_7�7g8989D9P9�9+:�:";�;K<=�=>�>�? � @   "0�01�1�1�2�4�4�4�4O6�6�7k8�8_9�9b:�:K;�;~<={=�=?E?�? � <   �021�1�24�4k6�6R7�7R8�8[9�9h:�:b;�;Q<�<X=�=O>�>�?   � @    000�0�12�4/5�5;6�6K7�728�8f9:�:N;�;O<�<?=�=?>�>;?   � @   �3�3�3�3�3�3�3�3�34<4H4#57(747[8�8�8"9'9�9:�:2;�;h<�< �    �2 7?>    P   �4�4l5{5�5�5�5�5�566%6c6k6}6�6�6�6�6�6�6�6 7�9_:�:2<�<�<_=�=>$>->�>     $   02X2d2O9�9s:;�;^<�<o=>�>�? 0 T   (0�0(1X2�2�3k4�4K5�5?6�6;7�7j8�8O9�9:�:�;<�<�<�<3=X=d=p=>>?>�>�> ??�?   @ L   0�01�112�233{3�3\4a4{4�4V5`5e5�67�78�9':�:K;�;K<�<?=�=?>�>B?�? P @   =0�0�1_23t3[4?5�526�78�8w9�9?:�:;o;�;L<�<+=�=J>�>4?�? ` H   0�01�1 2�2 3�34{4�4o5�5g6�6_7�7O8�849�9$:�:;"<;=�=>�>?�?   p L   0�01�12�23�34�4�4R5�5O67�7�7h8�8H9�9*:�:;x;�;x<�<x=�=x>�>x?�? � P   {0�0[1�1;2�23�3�3k4�4K5�5+6�67{7�7[8�8;9�92:�:;;{;�;�<R=3>X>d>�>O?�? � H   O0�0O1�1/2�2/3�3+4�4"5�56�6�6o7o8�8�8�8�8�8O9�9O:�:R;7<\<h<t<   � ,   �5�5�5�5�;�;�;<<#<f<v<�<�<�<�<�=P> �    �3�3q7�7�7@9Q9k9 � 8   h1m1~1�1�1�1'5�6Z8j8z8y9�9�9=:M:]:�<= =,=8=D=P= � 4   �1�1�1�2"5'585t5y5�5�5�5�5q7v7�7�7�7�7l=�=�= �     #1�1�1�1�1�1'4�4�6�6�6   �    p:�:h;�;(<�<      Y1^1v1a=�=�=?D?P?    �   O0J3w3�3-4j4�4�45B5u5�5�5'6p6�6�6(7r7�7�7888d8�8�8�8(9X9�9�9�9:H:x:�:�:&>+>2>9>@>G>N>U>\>c>j>q>x>>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>?Q?�?�?�?   T   0C0s0�0�07#7L788<8h8;9C9Q9�94:�;�;�;�;#<d<v<�<�<�<�<==+=�=�=�>?�?�?�? 0 h   V0e0�0111'1N1�12�23n3>4N4g4s4�455I5�6�6�678D8U8�9�9):i:�:;#;*;3;<;F;u;�;�;�;�;�;"=�=�>�>   @ h   ~23373?3�3�3�3F4U4w44�4�4�4�5�5�5�566-6�67.7�7�7�78#8N8�8�8,9x:}:�:�:(;-;�;�;�>�>?^?j?�? P ,   �5�5 6�67@768E8�8w9�9::%;3;i<6=�? ` $   �14(4�457�7�:u<6?H?�?�?   p     w26&898�8V9V:h:�:�?�?   � L   0F1U1j1q1�1�2y3�34v4�4�45*5{5�5�5/6y6�6�6/7H7�7�7�7H<�<=!=�>�>? � 8   �0�01V2e2�2�3�3'595w6�6�7�7�7�9�9�9&;5;Q;�<�<�< � @   �0�071Q1�1�2G3c3q3�3�3:5�6�6�6�67w8�8�89�9�9V:h:�:�>�> � (   �0�3�4G5�;�;�;"<R<�<�<4=�=>�>�> �     V2e2F5U568E8&;5;b>�>�?   � 0   j0	191'22�68f9u9�:�:�<�<�=�=�>�>�?�?   � �   F1U1w11�1�1�1�2�2�2�233-3�3�3�3�3F4S4m45575?5�5�5�5F6U6w66�6�6�6�7�7�7�788-8�8�8�8�8F9S9m9::7:?:�:�:�:F;U;w;;�;�;�;�<�<�<�<==-=�=�=�=�=F>S>m>??7???�?�?�? � �   F0U0w00�0�0�0�1�1�1�122-2�2�2�2�2F3S3m34474?4�4�4�4F5U5w55�5�5�5�6�6�6�677-7�7�7�7�7F8S8m89979?9�9�9�9F:U:w::�:�:�:�;�;�;�;<<-<�<�<�<�<F=S=m=>>7>?>�>�>�>F?U?w??�?�?�?     d   �0�0�0�011-1f2s2�233>3�3�34#4�4�4�5�5&959}9�9�9v:�:;;�;�;�<�<�<6=E=�=�=f>u>??�?�?�?  �   0#0N0�0�0�061C1n1�1�1�1V2c2�2�2�23v3�3�344>4�4�4�4&535^5�5�5�5c6�6�6#7F7S7~7�7�78f8s8�8�89.9�9�9�9:#:N:�:�:�:6;C;n;�;�;�;f<s<�<8=h=�=�=,>�?     t   0<0|0�01|1�1�12<2l2�2�2�2,3\3�3�3�34L4|4�4�45�5�6�<�<==h=m=�=�=N>S>`>m>r>{>�>�>�>N?S?`?m?r?{?�?�?�?   0 x   X0]0�0�0w1|1�1�1�1�1�1�1�1g2l2y2�2�2�2�2�2�2%3*3u3z3�4�4F5U5�5�5�6�667E7�7�7999 9%919M9R9W91:6:C:P:U:a:}:�:�: @ @   �7�7�7�7�7�7�7�7�7`8e8r88�8�8�8�8�8�8	9:!:&;9;;<Q<W=�= P     63H3b3�3�3/4:(:B:�:�:; ` L   �12@263E3�3v4�4�46%6`6�7�7 8�89@96:E:}:v;�;�;�<�< =�=>@>6?E?�?   p X   v0�0�0�1�1 2�23@364E4�4v5�5�5�6�6 7�78@869E9�9v:�:�:�;�; <�<=@=6>E>�>v?�?�?   � 0   �0�0 1�12@2�34(4;5I5�6i7":�;v>�>�?�?   �    �0�1�4N6�8�8�9�9<.= �    {0�2�5�5�6�69.:{=�? � $   �2�2�457(7�7�7�:�>�>[?i?   �    O2W6�8V;h;�;�<�<z=�= �     a4�4r7�:�:�:�:�:F?X?�?   �     �0�0j1q1Q8�8b;�>�>�>�>�> � $   �3;;�;�<�<F=V=>�>�>�?�?     <   �0W1�2�2�2�3�4�4,5�5�6�6j7�7�7J8�8�869E9f:x:�:�?�?�?  \   &585z5�5�516�6�6�6A7]7�788s8�8�839�9�9�9@:Y:�:�:;m;�;�;/<�<�<�<A=]=�=>>q>�>�>     d   �1�1�142M2�2�23a3�3�3!4s4�4�435O5�5�56c6�6�67m7�7�7/8K8�8�89a9�9�9!:q:�:�:1;M;>�>�>7?C? 0 (   �0�0f1u1f4r4&525�6�6�6}:�:�<�<   @ 0   �2�2�2�2�2�23 3$3(3,303�6�6�6}:�:�<�<   P 4   �2�2�2�2�2�23 3$3(3,3037<�<(=H=h=�=H>�>n?   ` (   0n0.1h2|3�3C4�5�6-7�7<#<�<�<   p <   00v1�163E3�4�4f6u6�6V8e8�8F:U:q:�;�;�;G=Y=�>�>�?�? � 8   61E1a13313�4�4�4&686W6�9�9�9�;�;�;�=�=�=&?5?Q? � 8   �0�0�1	2G3Y3�4�4�4f6u6�6�78!8�9�9�9&=5=�=�=%>�> � �   *0g0�0�0T1'2D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�5�56 6�6M7�8�89X9�9�:�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<>>.>P> �     �5�5�5�5=1=�=�=�>�>�>�> � @   �0�0�0 1�23�3�3f4u4�4�4�5�5606j8�89)9�:�:-<G<�<=�=�> � @   }0�0M1g133335)5C588s8�8f:u:�:�:�:�<�<==�>?N?g?z? � H   '1A1�1�1j2r3�3�3404O4�57:7H7w7�799�9�97:U:�:�:;�=>�>�>:?   � T   B0�0�0�0 11�2�3
44G4f4�5�5W6u67%7�7�7�7�:�:�:;;!;+;�<=!=7=I=Q=[=-?�?     0   0}0�12�2}3&454V46666g8y8w9�9�:�:=;W;     �4�5F9U9      �0�2�2U9V;h; 0 D   �7�7�8J9V:e:�;<�<�<�<�<&=3=M=�=�=>>f>s>�>&?5?W?_?�?�?�?   @ �   f0u0�0�0�0�01�1�1�1�1&232M2�2�233f3s3�3&454W4_4�4�4�4f5u5�5�5�5�56�6�678%8�8�8�8F9S9~9�9�9:f:s:�:;S;v;�;�;<<><�<�<=L=|=�=�=><>   P p   �0�0�0�0�0�0�0�0�0�1�1F2U2�2�2�3�3
444(4D4I4N4�7�7�7�7�7�7�7�7�78%8`8�9�9�9�:;@;6<E<�<v=�=�=�>�> ?�? ` (   0@061E1�1v2�2�47(7R7�8�8:9A9   p 4   0�0+3�6�6�6�6�66;F;�;�<�<�=�=j>�>�>V?h?�?�? � P   0^0�0�01\1u1�12)2z2�2�203|3�3�334O4�4�45�67F7U7�7�7�8�8�8\<c<c>j>   � 4   �4�4�4�4�4�4�4 55555L:c:�;�;F=U=??�?�? � \   0�0
2G2�2�2434$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5v7�7�7�7�>!?�?�?�?   � <    0�12�2�2�2�2j4�5�5#6268%8n8�8�8F:U:q:�:�:�:v<�<�< �     u4F6X6�9V:};�<�<
>�>�?   � $   �0�0Z2�2	4545�9�9:?4?�?   �    �3A4F4O4�4�5�59D:�: �    71�627T7]7"8E8N8l>y>      L31;�;�=  $   32�4�4	5�56g7�7�7Y8h8�;�;        \21:�:�< 0    �3�4�476}6�6+7:79   @     �0B1W3�:D;�;=]=}=>>   P    �2�2�2�2�:�:�:�:�?�? ` �   D0K0e0l0�0�0�0�0�011 1&1f1k1}12222�2�2333/343�3�3�3L4R4X4^4d4j4q4x44�4�4�4�4�4�4�4�4�4�4�4�4�4�455&5�5�5�5�5�5�5�5�5�5�5�5�5�56	666!6'616;6P6U6�6�6�6�6�6�6�6�6�6�6�67	777!7,71777A7s7�7�7�7z8x9,:9:W:e:r:,;9;F;Q;�<   p �   0+090�122#2+2024282a2�2�2�2�2�2�2�2�2�2�2333 3$3�3�3�3�3�3�3�3�34A4H4L4P4T4X4\4`4d4�4�4�4�4�4�7�78.83888�8�8�8�8�8�899 9J9O9T9:7:�;�;�;u=�=�=�=�=�=�=�=�=>5><>@>D>H>L>P>T>X>�>�>�>�>�>?%?@?G?L?P?T?u?�?�?�?�?�?�?�?�?�?�?   � l   >0D0H0L0P0h3�3�3�3(4X4|4�45\5�5�5�5,6�8�8�8�8(9-929::-:j:o:x:�:�:�:==-=�=�=�=F>T>g>�>�>�>�>�>*? � �   f0k0}0�0�0�0�0�0�0e1q1�1�1�1�1�12!2&2f3k3}3�3�3�3�3�3�3e4q4�4�4�4�4�45!5&5�6�6�6�6�6�6777:7?7D7�7�7�7:8?8H8r8w8|8�8�8$909d9i9r9�9�9�9�:�:;J;O;X;�;�;�;�;<4<@<t<y<�<�<�<�<)>.>7>a>f>k>�>�>�>�>�>�>f?k?}?�?�?�?�?�?�?   � �   ?0D0M0w0|0�0m1r1{1,313:3d3i3n3�3�3�3�3�3�3#4(414[4`4e4�4�4�4888m8r8{8�8�8�8v9{9�9�9�9�9:::O:T:]:�:�:�:�:�:�:;;#;�;�;�;h=t=�=�=�=�=�=>$>)>�?�?�? � �   :0?0H0r0w0|061?1K1T1b1k1y11�1�1�1�1�1�1�1;2L2[2�2�2�2�2�253V3f3�3�3�355-5p5u5~5�5�5�5�5�5�5!6&6+6R6�6�6�6
7[7�7�7�7�7�7�78+8>9�9�9�9�9�9�9f:k:p:w:;;6;Y;e;�;�;�;�;�;�;�;�;.<M<Y<i<u<�<�<===M=R=W=\=�=�?�?�? � �   0�0�0191>1g1�1
252W2�2�2�2(3�3�3�3�4�4�45�6�6�6�677<7A7a7f7�7�7�7�7�7�7�7X8d8m8�8�89M9|9�9�9:`:�:�:�:�:�:<<-<c<h<t<�<�<�<�<�<�=�=�=�=T>d>t>�>�>�>w?   � �   �0�0�0�0�0#1(141a1f1k1�1�1y2�2�2�2�3�3�3�34	4?4D4P4}4�4�4�4�4�4�4 55�5�6�6
777<7A7p7�7�7�7�8�8�8�8�8999�9�9�9&:+:=:Q:�:�:�:�:�:�:�:�:;$;*;7;�;�;�;<`<}<�<�<�=�=�=*>/>4>n?s??�?�?�?�?�?   � �   02070<0�0242e2�2�2�2�2333J3O3[3�3�3�3f4$8�8�8�8
999H9M9R9&:+:=:�:�:�:�:�:�:;;#;=;];�;�;�;�;�;�;�;H<M<Y<o<�<�<�<==4=�=�=�=�=>>>:>~>�>�>�>�>�>�>�>�>�>?/?9?>?J?d?u?�?   � �   �1�1�12	22"2'232I2U2^2c2l2x2�2�2�2�2�23'3~3�3�3�324=4F4N4W4_4e4k4s4y44�4�4�4�4�45$5q6�6�6�677+7X7]7b7x7�7�7�7�7�7�7�7�7�788]8b8n8�:�;�;�;�;<�<�<�<�>�>�>?? ?6?B?K?Q?Z?f?o?�?�?�?�?     �   0)0�0�0�0�0�0%1*1611�1�1�1�1Y2a2m2y2�2�2�2�2�2�2�2�2�2�2�2�2�23#3v3{3�3�3�3�3�3 44'4,484R4X4a4q4z4�4"6N6�6`8e8!9>9C9F;Z;><>  �   u0�0�0�0�0�0�0�0�0�0�0�01
111*1.1<1@1N1R1�1�1�1�1�12d2l2�2�2�2�2�2373[3|3�4�4�4�455�5�5�5�57�8�8�8�89C9�9�9�9_:g:�:�:�:�:1;o;�;�;�;�;�;i<>�>?B?M?_?�?�?�?   T   0D0Q0^0k0�0�0�0�0�011-1I1r1�1�1�1�2�2�2�2)303F3K3]3�4�45�5�5�5�8�8"9�<�< 0     01�3�5�5�56F7K7]7�78   @    62;2M2�7�748 P X   U1�1�152u2�2�253u3�3�354�4�4�4\5j5�5�56*6|6�6�6�7�7�7�7�7u8%;1;�<�<�<�<�<=:?�? ` �   31b1�3�3�344-4k4p4u4�4�4�4�4k5p5u5�5�5�5�5�6�6�6�6�8�8�8�8�8�899#9Y9^9g9�9�9�9�9�9�9:::q:�;�;�;�;�;�;�=�=�=�=�=>2>7><>>�>�>�>�>�>�?�?�? p �  00!0�0�0�011191>1C1y1~1�1�1�1�1�1�12-22272�2�3�3�3�3.444n4t4�4�4�45N5T5r5�5�5�5�5>6D6X6~6�6�6�6�6�67747^7d7�7�7�7�78868^8d8~8�8�8�89.949X9�9�9�9�9�9�9�9�9::::$:):3:9:F:K:U:[:i:n:x:~:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;
;;;';-;;;@;J;P;^;c;m;s;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<"<0<5<?<E<S<X<b<h<v<{<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====%=*=4=:=H=M=W=]=k=p=z=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>)>/>=>B>L>R>`>�?�?�?�?�?   � p   .040~0�0�0�0�0 11!1>1D1u1�1�1�1�2�3a4]8b8k8�8�8�8�8�8�8999�;�;�;<c<�<�<�<�<�<�<Y=^=j=�=�=�=>>�>? � �   �4555u5z55�6T7Y7^7�7�7�7:9?9K9x9}9�9�9�9�9:::\:a:m:�:�:�:�:�:�:(;-;2;q;�;�;�;�;�;h<r<:>A>}>�>�>�>�>�>-?2?>?k?p?u?�?�?�?   �    $0)0.0�0�0�0�0�0�0s2x2�2�2�2�23$303]3b3g3�3�3�3444�4�4�4�4�4�4M5R5^5�5�5�56
66C6H6M6�6�6�6�6�6�6�7�7�7�7�7�7:8?8K8x8}8�8�8�8�8999�9�9�9�9�9�9.:3:?:l:q:v:�;�;�;�;�;�;t<y<�<�<�<�<K=P=U=>>>8><>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>   � L   w58#8B8�8�9�9�;�;�;�;�;�;�;�;�;�;�;(<,<0<4<8<<<@<D<�> ??
?p?u?z?   � �   1p1u1z1�1�1�1b3444�4�4�4j5o5t56"6'6�6�6�6r7w7|7 88
8�8�8�8f9k9p9,:1:6:�:�:�:�;�;�;~<�<�<$=)=.=�=�=�=N>S>X>�>�>�>   � H   �2�2�2 3%3*3p3u3�3�3�3�3444D4I4N4�4�4�4(5-525W6\6h6�6�6�66;8? � h   �0�0�0�0�0�2�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8:�:�:;;g<
=0=�=   � �   30�0>1D1�12O2T2Y2�23G3M3m3t3z3�3�3�34>4D4}4�4�4�4.545T5�5�5�5�5�536�8�8�8�8F9K9]9�9*:9:X:e:s:�:�:�:�:�:�:�:�:�:�:;;+;B;p;<<0<z<�<�<=F=�=�=j>�>�>?F?�?�?�?�?   �    0�0�0"1S1�122.2T2]2c2�2�2�2�2�2�2�2333r3�3�3
4\4�4�4�5�5�5666"6,6h6x6}6�6�6�6�6�6�64797>7C7M7j7o7t7�7�7�7�8-9j9�9	:::�:w<�<�<�<�<�<�<1=6=B=o=t=y=�=�=�=�='>1>??!?N?S?X?�?�?�?�?�?�?�?    �   (070N0�0�0[1c1l1v1�1�1�1�12+252j2y2�2�2�2�2�2�2�2�2�23'3:3Q3Z3j3n3x3�3�3�4�4�4�4�4�4�4�4�4�45�5�5�5�5�566=6B6N6{6�6�6�677*7W7\7a7y7�7�7�7�7�7�7�7X8�9�9�9�9�9�9�9�9::b:�:�:�:�:�:�:�:�:�:�:K;�<z=�=�=�=	>�>   8   �2�2�3M425A546?6e6p6�6�6�6�6a7E9�9p>?�?�?�?�?   0 �   �2�2f3�3�3�3�3�3
4Z45�5�5�5W6d6m6u6�6�6�6�7�7>8F8d8m8u8�8�8�8�8�8�8�:�:�:;;;T;\;�;�;�;�;�;�;r<z<�<�<�<�<===P=W=�>�>�>�>�>�>??-?v?�?�?�?�?�?�?   @ �   070<0E0z00�0�0�0�012&2\2o2�2
333�3�3�34.434<4f4k4p4�4�4�4�4�4�45<5Y5c5�5�5�5�6�6�6�6	777L7Q7V7|7�7�7�7�7�7�7-8v8{8�8n9�9�9�9.:3:8:^:�:�:�:;;;6;|;�;�;(<�<�<�<==4=n=>2>?Y?c?�?�?�?   P `   70�01+1^2h2�2�3�3	4&5;5�5�5�56$6F6�6�:�:�:�:�:�:A<M<�=�=�=�=�=>>4>�>'?:?W?l?r?{?�?   ` X   l0�0�0K1h1�12�3�3�3	44*4v4{4�4�4�4�4	555�5�5�5�5�677�7�7T8^8l9�9�:\<�>�>�>   p �   Z0_0k0�0�0V2[2m2�2�2�2�2&3+303Y3�3�3�3�3�3�34d4i4r4�5�5�5�5�5�56m6r6{6�6�6�6f7k7}7�7�7�7�78(838H8�89979<9A9�9�9�9�9�9:::�:�:�:;;;?;D;I;�;�;]>b>n>�>�>�>�>�>�>??$?   �    �1�1222!262;2M2�2�2�2�2�2v3{3�3�3�3�3414N4�4�4�45
55)5�5�5�5�5l6p6t6x6|6�6�7�7�7�7�7w8�8�8�8�8�8�8�8�8�8�8999#9+929E9J9R9Y9l9q9�9�9�9:	:l:�:�:�:�:�:;;;D;H;L;P;T;p;t;�<�<�<�<�<�<�<�<==6=;=@=J=Q=V=[=e=l=q=v=�=�=�=�=�=�=�=�=�=�=�=�=8>B>`>y>�>�>�>�>�>�>
??+?6?=?U?\?   � �   �0�011A1F1K1j1v1�1�1�1�1�12!2o2t2}2�2�2�2�2�230353:3W3c3s3�3�3�3�4�4�4�455.5;5@5F5S5X5^5�5�5�566$6)6\6h6t6y6~6�6�6�6�6�677757:7?7D7�7�7�7�7888$8O8T8Y8�8�8�8�8�899+949f9�9q:�:�:�:;;;);3;};�;�;<f>k>�>Q?o?t?y?�?�?�?�?�?�?�?�?�? � �   d0i0n0�0�0�0�0�0�0�01181=1B1v1�1�1�1�1�1�1�1�1+2_2d2i2�2�2�2�2�2�2�23"3'3n3s3x3}3�3�3�3P4�4	5=5P5a5h5�5�5�5�5�5�5X6_6�6�6�6�6�6777�7;�;C=�=C>H>T> � �   10111G1h1[2�2�2�2�233&363D3H3L3P3T3�3�3�3�3�3 4*4O4�5�5
6#66:;:M:w:�:�:�:�:&<+<=<�<�<==b=n=}=�=�=>>$>(>1>C>w>g?�? � �   0�01H1b1�2�3�3�3B4G4P45!5,737B7�7�788D8�8�8�8999X9_9q9x9�9):0:;;-;p;u;~;�;�;�;�;�;�;!<&<+<R<�<�<�<
=[=�=�=�=�=�=�=>+>>?�?�?�?�?�?�?   � �   d0i0n0v0�0	111T1`1}1�1�1�1�1�1�1�1)2H2T2d2p2�2�2333H3M3R3W3~355%565;5M5,6s6�6�6�7�7�788@8^8�8�8�899-9F9�9:�:�:�:�:	;3;�;�;�;�;�;�;�;�;?<F<S<X<�<�<�<�<�<6=v=}=�=U>]>b>k>�>�>�>�>�>V?[?m?�?�? � �   000�0�0�0�0�013181�1�12333�344#465;5M5�5�5�5�5�5�6�6�6�6�6#7(747�7�7�7�8�8#;(;4;a;f;k;�;�;�;�;�;<_<d<p<�<�<�< � h   l5q5}5�5�5�5�5�5686=6B6�6�6�6�6�6�6�7�7�78�8G:�:�:�:�:�:�:#;(;4;a;f;k;q=v=�=�=�=�=�=>>=>B>G>   l   w0�0�0�0111S1X1d1�1�1�1'3�3�3�3�3�3�3444E4J4O4::":�:�:�:O;c;i;=�=�=�=>)>1>6>D>L>Y>e>�>??  �   �3�3J4i4o4�4�4�4�4555J5Y5l5�5666%6:6F6V6�6�67u7�7�7�7�7B8I8]8r8y8�89"9+9U9Z9_9�9�9�9�9�9�9I;�;X<�<>??-?5?E?V?   �   f0k0}0�0�0�0�0�0$141t1�1�1�1k2p2u2�2�2�3�3�34M4R4W4�4�4�4�4�4 5:6m6�6�6�6�6�6�6�6�6 77�7�7:8�8�8�89 9%9*9�9�9�9�:�:�:;@;E;J;�;�;�;�;�;�;<<<m<r<w<�<�<�<f>k>}>�>8?�?�?�?   0 d   0\1�1�132�3�3�3&4+4=4�4�4�4�4�4�45�5�5�56V7�7�7�7�7�7�7�8�8�89�9�95:A:�;�<&=@=i=�=�=�=   @ P   :12�2�2�2q4�4�5686D6�8�8�8�8�8�89�9�97;<;E;o;t;y;H<p<m=>�?�?�?�?�?�? P x   0#0�0�0�0�0�0�0h1p122\2a2m2�2�2�2�3�3*5w5|5�5�5�5�5�6}7�78�9�;�;�;�;�;�;9<A<�<�<�<�<�<=d=k=�=�=D>I>U>�>�>�> ` �   00-0o0}0�0�0�01161J1b1~1�1�1�1�2333*3/383S3X3a34	44<4A4F4�4�4S6X6d6�6�6�6�6777I7N7S7�7�7�7�7�7�7.8^8�8�8�8�899!9q9v9�9�9�9�9�9�9D:H:L:P:T:X:\:`:d:h:l:p:t:�<�<�=�>�>�>�>?	??�?   p �   "0�0�061@1"2�23�4�6�67J7O7X7�7�7�768;8M8�8�8�8�8�899,9W9\9e9�9�9�9�9&:+:4:;;@;I;�;�;�;�;�; <><�<�<�<�<�<�<=#=(=1=�=�=�=>>>t>{>   � |   $0)050b0g0l0�0�0�0�011$1�1�1�1�1�1�1�1/2_2�2�2�2�2�2�2B3G3S3�3�3�3�3�3444 4$4(4,4044484<4@4D4
:?:?}?�?�?�?�?�? � �   p0�0�0=1B1K1u1z11�1�1�1�1�1�1i3�3]4b4k4�4�4�4�4�4�4555�6�6757:7?7�7�7�7�7�7�78[8c8�8J9Q9�9�9�9�9�9�9':/:�;�;`<e<q<�<�<�<�<�<�<#=(=-=V=�=�=�=�=>.>3>8>v>~>�?   � t   S0X0d0�0�0�0$161x1�1�1�1�1222y2~2�2�2�2�23�3�3{4�4�4�4�4�4�5�5�6�6L8S8K9P:�:�;�;�;�;�;�;�<�=�=�=�= >'>   � h   054585<5@5D5H5L5P5T5X5\5`5d5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5h>�>�>�>�>�>�>???I?N?S?   �    �0�0�0111]1b1k1�1�1�1�3�3�3�3�3�34f4k4}4%5*5/5]5k5w5�5�5�5�5�5�5�5�5�5�5�5�5�56&61696A6I6S6[6c6�6�6�6�6�6�6Z7`7n7|7�7�7�7�7�7�7"8-8G8�9�9�9&:+:=:�:�:�:�:�:�:�:�:;%;/;8;=;B;g;q;�;�;�;�;�;�;�;�;�;�;�;<+<�<�<�<�<==0=O=U=m=r=w=�=�=�=�=]?b?g?   � �   �1�1{2�2�2�23-353C3_3k3p3u3�3�3�3�3�3�3�3�3�3�3�3�3�4�4�4�455'5Q5V5[5r5�5�5�566626�6�6�6�6�6�6�6k7p7y7�7�7�7�7 8	83888=8|8�8�8�8�8�8�89:?E?^?r?x?~?�?�?�? � �   00�0�0�0�0�01#151G1d1z1�1�1<2H2T2`2l2x2�2�2�2�2�3�3�3�4�465?5L5V5^5c5j5�5�6�6778$8-8W8\8a8�8�8�89959:9?9�9�9�9:: :J:O:T:�:�:;0;5;>;h;m;r;�;�;H=M=V=�=�=�=�=�=5><>�>�>�>�>�>�>F?K?T?   � �   00<0e0j0s0�0�0�0�0�0G2y2�2�2�2�2�2�2�2�2�3�3�3�3�3�3	44o4w4�4�4�4�455}5�5�556=6h6�6�6�6�6�6�677L9o9�:�:�:;�<�<�<=='=Q=V=[=�=�=�=�=�=�=�=�=> >%><>F>x>}>�>�>�>�>�>�>�>�> ??�?�?     �   0�0�0�0&1.1M1W1v1�1v2{2�2�293D3�3�3�3'484P4�4�4)5R5z5�5�5�5�577C7O7v7�7�7�7E8h8m8y8�8�8�8�8999U9Z9_9�9�9�9:o:~:;1;N;h;�;�;�;�<�<�<== =6=�=�=�=>!>*>T>Y>^>�>%?*?3?  �   0�0�1�1�1f2t2�2�2�2�2�263Y3^3g3�3�3�3�3�3�34:4?4D4~4�4�4�4�4�45M5R5[5�6�6�6�67!7&7L7w7|7�7�7�7�78	88M8R8W8�8�8�8�8999D9�9�9�9�9�9�9!:~:�:�:�:�:;;B;f;�;�;�;-<o<�<�<=D=m=w=�=�=�=>>1>�>�>?'?E?�?�?�?     `   �0�0�0�0=1�1/2~2�2�23x3�3�3/4M4!5?5[5y5�5�5�5�6�6�687�7�7�7n=�=�=�=> >%>�>�>0?�?�?�?   0 �   000L0Q0]0�0�0�0�2�2�2�2�2�2%3*363c3h3m3�3�3�3i4�4�4@5E5Q5~5�5�5�5�597�7-828>8k8p8u8�8�8�8�8�8�8	;k;�;�;�;<#<(<e<j<v<�<�<�<�<=!=t=y=�=�=�=�=�=>?�?�?�? @ L   000|0�0�0�0�0�0�1�1�1�2�2�3�3N5U5�6�7!8�8�8�8,91969?:�:�:5;<;|;�; P �   �2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 3$3(3,3034383<3@3D3H3L3P3T3X3�:�:�:�:�:�:$;,;y;~;�;�;�;�;.<5<`<�<�<�<�<�<�<F=M=x=�=�=�=�=�=�=#>+>�?�?�?�?�?�? ` �    0%010^0c0h0�0�0111K1P1U1�1�1�1�1�1�1�2�232373<3Y6^6g6�6�6�6�6�6�6777O7V7�7�7�7�7�7�7<8A8J8t8y8~8j9o9{9�9�9�9?;D;P;};�;�;�;�;�;�;<<C<K<�<�<�<�<�<�<9=>=J=w=|=�=�>�>�>�>�>�> p t   	222A2F2K2�2�2�2�2�2�23	3p3u3~3�3�3�3�3�3�3)4.434(5-595f5k5p5�6747S7r7�7�7�7�78,8K8j8=9e9�9-=�=�=�=�=   � ,   �0�0�0�01�1�1E2�3�3�3�3�3�344+4   �    �1.2;2m2r2{2 �    �566�6�6�6<   � l   1�2|4�4>5D5J5Y5a5i5s5�5�5�5�5�5�566�677�7�9{=�=�=�=�=�=�=�=8>E>K>p>�>�>�>?#?6?=?B?W?]?j?p??�?   �    �3y4B5d6"808b8+=_=   �     �2�2�4x5�5�5�8:;<�=.? � 0   H192Q3^4$5O5�<�<�<=5=e=�=�=�=%>T>t>�>P? �    %0U0�0�0�01f1x1�1�1�1�1�1�12#262M2�2 3	33"3<3E3J3{3�3�3�3�3�3�3�45F5@6j7w7�7�7�7�7G8X8c8l8�8�8�8�8�8�8�8	9989J9S9m9t9�9�9�9�9�9�9�9:::l:�:�:�:�:�:�:);0;9;Y;�;�;�;<<n<�<�<�<�<�<�<�<�<�<�<�< ==(=,=0=4=8=<=@=D=H=L=P=T=X=�=�=�=�=�=�=�?�?�?�?�?   �   0�0�0�0�0�0�0 111�1�1�12�3�3�3�34#404945-5�5�5�5�5�5x6�6i:�: ;	;;5;L;U;\; <*<><J<i<z<�<�<�<�<�<�<2=C=r=|=�=�=�=_>l>z>�>�>�>    �   0!0'00050Y0k0�0�0�0�0�0�0*1<1]1j1�1�1�1�1�1�1e3r3�3�3�3�3�3�3�3�3�3x4�4�4�4�4�4�4�4�4�4�45555�5�5�5�5�5�5�5�5�6�6�6�6�67717=7F7e7l7u7�7�7�7�7�7�7�7�7�7�7O8W8]8�8�8�8�8�8�8999'9<9|9�9�9�9 :::4:A:J:);�;<<,<L<Z<b<n<z<�<�<=4=�=�=�=�=?   �   �1�3�4�4�4�4�4�455-5:5M5c5k5s5~5�566676>6C6K6�6�6�6�6%7>7�7�7�7�7�7�788%8+848T8_8z8�8�8�8�89&9D9O9�9�9�9:I:X:c:k:�:�;�;�;�;<<'<@<H<a<�<�<�<�<�<�<�<=&=5=[=i=r=�=>4>8><>@>D>H>L>�>�>�>�>�>�>�>�>�>�>�>�>�>D?H?L?P?T?X?\? 0 �   �12_2y2�2�2�2�2�23'3c3l3r3�3�3�3�3�3�3�3�3�314`4h4o4�4�4�4�4�455 5$5(5p5t5x5|5�5�5�5�5�5�6�6�67717K7X7`7�7�7g8x8�8�8g:x:�:�:�:�:�:�:;,;W;<<<�<�<�<�<�<&=8=A=F=i=p=}=�=�=�=�=�=�=D>M>�>�>�>�>�>�>,?5?j?�?�? @ �   0w0�0111111�2�2�23 3)303h3�34#4,4,5�5D7O7W7c7n7v7�7�7�7�7�7�7�7�7�788�8�89!9�9�9�9�9�9:::4:I:W:e:x:�:�:�:�:�:�:�:�:�:�:�:;%;g;�;�;�;�;<<&<b<u<j=t==�=�=�=�=�=�=�=>�?�?�? P �   00�0{1�1�1�1�1�1�1�1�1�1�1�14282<2@2D2�3�3�3�3�3�3�3%404<4V4d4m4�45 5(515:5B5�5'646B6K6{6�6�677%767H7W7`7�8T9i9q9w9�9�9::#:):2:8:R:Y:^:f:v::�:�:�:�:�:�:�:!;);8;A;G;U;b;�;�<===0=;=C=r=�?�?�?�?   ` �   0000000 0$0(0,0004080<0@0D0�0�0�0�0�01111111 1$1�3�3�3�3s4�4�4�45f5w5�5�5�5�5�56666W6e6n6'717H7Q7_77�7�7�7�7�7�7888!8*83898M8R8Z8�8�8�8�89C9b9k9t9�9�9�:>>#>.>7>E>Q>]>i>�>�> p \   f1k1}1�1 2v2{2�2�23�3H5M5V5�5�5�5�5�5�5�5 66g6l6u6�6�6�6�6�6�677$7�8g:<?v?{?�? � d   2'2S2X2a2�2�2�2�2;3@3I3s3x3}3=4�4�5�5�5�5 66666�8�8�8�8�9�:�;�<�<�<}=�=�=�=>>6?;?@?   � L    00
0}0�0�0Z2�2�2�2�3&4/4�4�6�677�7�7�7�7�9D:�;�;�;�<�<�=�=�>?�? � D    1J4�4U7}7�7�7�7A8�8�9�:�:�:;�;�;Z<<v={=�=�=�=�=>>!>�>�> � x   000a0f0r0�0�0�0�0�0�0)1.131{1�1�1�1�1�172Y2�4�4�4�4�4�4"5'505Z5_5d5�8�8�8�8�8�8C9H9Q9{9�9�9�>�>�>�>S?�?�?�?�? � �   0070<0A0�0�0&2+2=2�2�2�2�2�2�2333I3N3S3�3�3�3�3�3�3W4y4�5�5�5�6�6�6�6�6 71787�7�7�7888999O9T9Y9�9	;+;5;i;�;�;�;�;<<*<�<�<�<V>[>g>�? � �   20111�1�1�1D3m3�3�3 4"4Q4�4�4�45,5054585<5@5�5�5�5�5�5�5�5�5�5�58:w:|:�:�:�:�:�:�: ;*;/;4;�<�<�<===E=J=S=}=�=�=�? � �   �0�0�0�0�0�0~1�1�1�1*2/2;2k2p2u2�2�2�2333p4�4�5�5�56
66�6�6�6�6�6�6J7888L8Q8V8!9(9::?:K:{:�:�:�;�;�;�;�;�;G=L=X=�=�=�=�>�>�>�>�>�>�?�?   � �   !1(1�1�1�1222�233=3B3G3F4K4W4�4�4�4|5�5�5�5�5�5�6�6�6�6�6�6�7�7�7+80858�8�9�9�9:$:):;;%;U;Z;_;�;[<(=-=9=i=n=s=^>c>o>�>�>�>D?I?U?�?�?�?     �   {0�0�0�0�0�0�1�1�1�1�1�1�2Q3V3b3�3�3�3�3�3�3u4|4�4�4 55�6�6�6�6�6�6�7�7�7888�8�891969;9&:+:7:g:l:q:^;c;o;�;�;�;�<�<�<�<�<�<�=�=�=�=�=�=�>�>�>)?.?3?  �   00%0U0Z0_0J1O1[1�1�1�1e2j2v2�2�2�2�3�3�3�3�3�3�9�9�9�9�9�9~:�;�;�;�; <<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=h=l=p=t=x=|=�=�=   0 t   �2�3�3�3�3�3�3t4�4�4�4 5%515a5f5k5�5�5�5
666�67O7T7`7�7�7�7�7�8�8�8�8�8�8�9�9�:�:Q<X<P=U>�>�?�?�?�?�?�?   @ h   �0�1�1�1�1%2,2G9L9X9�9�9�9�9�9�9�9�9�9 ::::::::4:8:<:@:D:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:   P T   �2�2�3 4$4;4f4k4}4�4�4�4�4�4�4M7R7[7�7�7�7L8Q8Z8�8�8�8949�9�9�9�9�9�96?;?M? ` �   00*0W0\0a0�0�0�0�0�0�0�1�1�1G2P2f2233*3�3�3�344!4u4z4�4�4�4�4/54595�5�5�5*6/686b6g6l6�6�6�6�6�6�6�7�7�7�89o9t9}9�9�9�9�;�;<<D<q<�<�<�<�<�<�<-?5? p �   -050A1H1�1�12 2}2�2�2�283=3I3v3{3�3�3�3�3�3 44�5�5�5�56	66�9�:�:�:;#;(;�;�;�;�;�;�;%=[=y>~>�>�>�>�>f?k?w?�?�?�?�?   � �   �0�0�1�1�1/24292M3R3^3�3�3�3�455>5C5H5\6a6m6�6�6�6i7p7�8�8k9p9|9�9�9�9�:�:�:�:�:�:r<w<�<�<�<�<�=�=�=�=�=�=j>�?�?�?�?�?�?   � �   �0�0�0111�152333O3T3Y3F4K4W4�4�4�4,515=5m5r5w5d6i6u6�6�6�6�7�7�7�7�7�78<9A9M9}9�9�9�9�9�9`:g:�:�:�:�:�<�<�<�<�<�<�=�=�=�= >>�>�>�>%?*?/? � �   0!0-0]0b0g0T1Y1e1�1�1�1�2�2�2�2�2�2�3�3�3�3�3�3�4�4�4#5(5-5666O6T6Y6F7K7W7�7�7�7a8f8r8�8�8�8�9�9�9�9�9�9�?�?�?�?�?�? � h   {0�1�1�1�1�1�1<2@2D2H2L2P2T2X2\2`2d2h2l2p2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33@3D3H3L3P3T3X3 � T   �3C4H4T4�4�4�4�4�4�4-52575�5*6t6y6�6�6�6�67�7�799s:z:�;�<F=>>!>Q>V>[>d? � d   00Z0a0�0�0�7�7�7	888h8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,909 � 4   �011r1~1D2P2V4[4m4�4�4�4�4�4�4�:D>d>�>�?   � ,   W0g5q5�5�7q8v88�8�8�8H9a:h:�;�;�<�<   X   �1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1222L2P2T2Z5�6�6�6�67777b7g7l7q7�7�7�7�7    D   �0�5�6�6�6�9�9�9�9<:�;H>v>{>�>�>�>�>�>�>?5?:???{?�?�?�?�?�?   �   �0�0�0�0�01G1L1U11�1�1�1�1�1
222�4�4�5�56V6V7[7m7�7�7�7�7888E8p8u8~8�8�8�8�899A9F9K9�9�9�9�9�:�:
;7;<;A;X;�;�;�;<<<-<v<{<�<�<�<�<)=.=3=k=�=�=�=�=�=�=�=!>&>/>Y>^>c>�>�>�>�>�?   0 �   0�0�0�0�01(1G1h1�1�1�1�1�12�2�2I3N3W3�3�3�3�3�3�34!4&4u9�9�9�9@:n:�:�:�:&;+;=;�;�;�;�;�;�;�<�<�<K=P=Y=�=�=�=�=�=�=(>->2> @ T   �3�3�4�4�6�6�6;7R8W8`8�8�8�8�8�8�8999e9j9s9�9�9�9W;\;e;�;�;�;�;�;�;<<< P H   �0�0�00252A2�2�2G4�56[6`6i6�6�6�6 77787=7B7�<�<�<==�=�=�>? ` �   '1s1x1�1�1�1�1�2�2444@4E4J4�4�4�4�4�4�4/555=5K5Q5d5�5�5�5�5�5�5�5�566!63686D6�6�6	7`7q7�7�7 8%8*8�8x:�:�:;;�;�;<E<�<�<�<==$=j=o=x=�=�=�=�=�=>->2>7>   p D   �3#4(414[4`4e45$5'6�7�7�7�7�7�7W9b:�;z<1=6=?=l=q=v=
>$?+?   � �   y0�0c1j1\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6 7$7(7&:,:2:8:>:D:J:P:V:\:b:h:n:t:z:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;
;;;;";(;.;4;:;@;F;L;R;X;^;d;j;p;v;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<$<*<0< � �   �2%3U3�3�3454o4�4�45*5I5l5�5�5�56=6�6�6�67J7z7�7868v8�8�89V9�95:�:�:/;j;�;�;�;�;<#<J<�<�<$=d=�=�=$>�>�>"?d?�?�?   � �   $0�0�0C1�1�1�12J2z2�2�2
3:3j3�3�3�3*4Z4�4�4�45J5z5�5�5
6:6j6�6�6�6*7Z7�7�7�78J8z8�8�8
9:9j9�9�9�9*:Z:�:�:�:;J;z;�;�;
<:<j<�<�<�<*=e=�=�=
>:>j>�>�>�>"?�?�?   � �   &0f0�0�01i1�1�1&2f2�2�23C3c3�3�3464v4�4�45V5�5�5�566f6�6�67F7�7�7�7&8f8�8�89F9v9�9�9&:V:�:�:;6;v;�;U<�<5=z=�=�=?>�?   � �   �1\2�2�2�223b3�3�344�4�4�4�45'5B5]5x5�5�5�5�56�6�6�6�6�67"7=7X7s7�7�7�7�7�8�8�8*9�9�:d;�;�;$<d<�<�<$=d=�=�=P>�>�>?T?�?�?     �   0�0�0�01J1z1�1�1
2L2�2�2<3�3�3,4|4�4$5u5�5�67Z7�7�7�78J8z8�8�8
9:9j9�9�9�95:j:�:�:�:I;s;�;�;<F<�<�<�<&=f=�=�=>F>�>  P   0�0�0
1#1;1S1k1�1�1�1�1�1b2�2h3�34J4z4�4�45l5�56�6�67J7a7i7�7�7�78   L   ;o;�;<_<�<�<�<�<=4=T=t=�=�=�=�=>4>T>t>�>�>�>�>?4?T?t?�?�?�?�?   0    040T0t0�0�0�0   P �   111111 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�2�2�2�2�2�2�2�3�3�3�3�3�3�3�3�3�3�3�3 4444444 4$4,40484<4D4H4P4T4\4`4d4l4p4x4|4�4�4�4�4�7�7�7�7�:�:�;   ` $  (0,0004080<0@0D0H0L0D1H1L1h1l1p1t1|1�1�1�1�1�1�1�1�1�1 2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�233333 3$3034383D3H3L3T3X3\3`3d3h3l3�3�3�3�3�3�3�3�3�3�3�3�3�3�34444 4�4�4�4�4�4 55555555 5$5(5,5054585H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�8�8�8�8�8�8�8�8�8�8�8 p �   t3x3H4L4P4X4\4d4h4l6p6x6|6�6�6�6�6�7�7�7�7�7�7�7�7�7888(848@899 9,989D9P9\9h9t9�9�9�9�9�9(<,<0<L<P<T<\<`<d<l<p<t<|<�<�<�<�<�<�<�<�<�<�<�<   � @  �3�3�3�3D4L4T4\4d4l4t4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�45555$5,545<5D5L5T5\5d5l5t5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56666$6,646<6D6L6T6\6d6l6t6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67777$7,747<7D7L7T7\7d7l7t7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78888$8,848<8D8L8T8\8d8l8t8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89 � x  44 4$4(4,4044484<4@4D4H4L4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�6�6�6�6�6�6�6�6�6�6�6�6�6�6�677777 7$7(7,7074787H7L7P7T7X7\7`7d7h7�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>> >$>(>,>0>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>?? ?$?(?,?0?4?8?<?@?D?H?L?P?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   � t   000000 0$0,0004080<0@0H0L0P0T0X0\0`0d0h0l0p0t0x0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0111111 1$1(1,101<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 222222 2$2(24282<2@2D2H2T2X2\2`2d2h2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3034383<3@3D3H3L3P3T3X3d3h3l3p3t3   � �   �0�0�0�0�0�0�01111111(1,1014181<1D1H1L1P1T1X1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222 2$2(2,2024282<2@2D2H2T2X2\2`2d2�8�8�9�9�9�9�9�9�9�9 ::::   �    44 4P<T<X<\<`< �    �1�1�13333     �  X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5(50585@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6h6p6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 8888 8(80888@8H8P8X8`8h8p8x8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 9999 9(90989@9H9P9X9`9h9p9x9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::: :(:0:8:@:H:P:X:`:h:p:x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;`;h;p;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<<$<,<4<<<D<L<T<\<d<l<t<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====$=,=4=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   0 �   0000$0,040<0D0L0T0\0d0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01111$1,141<1D1L1T1\1d1l1t1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222$2,242<2D2L2T2\2d2l2t2|2�2�2�2   @ L    1$1(1,1014188888,:4:<:D:L:T:\:d:l:t:|:�:�:�:�:�:�:�:�:�:�:�:�: p    �=�=�=�=@?D?H?   � ,   80@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0   � �   �5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7   � �   22 2$2,2024282@2D2H2L2T2X2\2`2h2l2p2t2|2�2�2�2h6t6�6�6�6�6�6�6�6�6�6�6�6777(747@7L7X7d7p7|7�7�7�7�7�7�7�7�7�7�7 888$808<8H8T8`8l8x8�8�8�8�8�8�8�8�8�8�8�899 9,989D9P9\9h9   � 8   03<3H3T3`3l3x3�3�3�3�3�3�3�3�3�3�3�344 4,484    (   t5,?D?\?d?x?|?�?�?�?�?�?�?�?�?     �   000,04080@0X0d0|0�0�0�0�0�0�0�0�0�0�0114181L1T1\1t1�1�1�1�1�1�1�1�1�1�1�12 2,2D2\2`2t2|2�2�2�2�2�2�2�2�2�2�2�2�23$3(3<3D3H3P3h3�3�3�3�3�3�3�3�3�3444 44484L4T4X4\4d4|4�4�4�4�4�4�4�4�4�4�45555 5(5@5X5\5p5x5�5�5�5�5�5�5�5�5�5�566(6064686<6D6\6t6x6�6�6�6�6�6�6�6�6�6�6�6 770747H7P7T7X7`7x7�7�7�7�7�7�7�7�7�7�7�7 888 8$8(808H8`8d8x8�8�8�8�8�8�8�8�8�8�8�8 990949H9P9X9p9�9�9�9�9�9�9�9�9�9�9::$:<:@:T:\:d:|:�:�:�:�:�:�:�:�:;;;;0;H;L;`;h;l;t;�;�;�;�;�;�;�;�; <<< <$<(<0<H<`<d<x<�<�<�<�<�<�<�<�<�<�<�<�<= =$=8=@=D=H=P=h=�=�=�=�=�=�=�=�=�=�=�= >>>$><>@>T>\>`>d>l>�>�>�>�>�>�>�>�>�>�> ??? ?$?,?D?\?`?t?|?�?�?�?�?�?�?�?�?�?�?�?�?   0 �  0 0$080@0D0H0L0T0l0�0�0�0�0�0�0�0�0�0�0�0 11111141L1P1d1l1p1t1|1�1�1�1�1�1�1�1�1�122$2,20242<2T2l2p2�2�2�2�2�2�2�2�2�2�2�2�2�23,303D3L3P3T3\3t3�3�3�3�3�3�3�3�3�3�34444444L4P4d4l4p4t4x4�4�4�4�4�4�4�4�4�4�455(5054585@5X5p5t5�5�5�5�5�5�5�5�5�5�5 66666(6,6@6H6L6P6T6X6d6|6�6�6�6�6�6�6�6�6�6�6�6777 7(7@7X7\7p7t7�7�7�7�7�7�7�7�7�7�7�7�7 880848H8P8T8X8`8x8�8�8�8�8�8�8�8�8�8�8�89999$9<9T9X9l9t9x9|9�9�9�9�9�9�9�9�9�9�9�9::,:D:L:P:T:X:l:p:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;$;<;@;T;\;`;d;l;�;�;�;�;�;�;�;�;�;�;�;<<,<4<8<<<@<H<`<x<|<�<�<�<�<�<�<�<�<�<�<�< == =8=<=P=X=\=`=d=h=t=�=�=�=�=�=�=�=�=�=�=>>>>> >,>D>\>`>t>|>�>�>�>�>�>�>�>�>�>�>�>�>? ?$?8?<?P?T?h?p?t?|?�?�?�?�?�?�?�?�?   @ P  00 0(0,00080P0h0l0�0�0�0�0�0�0�0�0�0�011 141<1D1\1t1x1�1�1�1�1�1�1�1�1�1�1�12,202D2L2P2X2p2�2�2�2�2�2�2�2�2�2�2333(366 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :,<<<h<p<�<�<�<�<�< =(=L=X=`=�=�=�=�=�=>> >H>l>x>�>�>�>�>�>?,?8?@?`?h?t?x?�?�?�?�?�?�?�?�?�?�?�?�? P �  00(040H0T0\0h0l0x0�0�0�0�0�0�0�0�0�0�0�0�011$181D1L1X1\1`1l1�1�1�1�1�1�1�1�1�1�1�1�1�1�122$20242@2T2`2h2t2x2|2�2�2�2�2�2�23383D3h3t3�3�3�3�3�3�344@4H4T4�4�4�4�4�4�4�4�4�4555(5P5\5�5�5�5�5�5�5�5�56646@6d6p6�6�6�6�6�6 7$7,787`7h7p7x7�7�7�7�7�7�7�78(80888D8l8x8�8�8�8�8�8�8�8�8$9,949<9H9p9|9�9�9�9�9�9�9:@:L:T:t:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;t;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<<H<l<t<|<�<�<�<�<�<�<�<$=0=T=\=d=p=�=�=�=�=�=�=>><>H>l>x>�>�>�>�>�>?,?8?\?h?�?�?�?�?�?�?�?�?�?�?�?   ` �  0$0P0X0|0�0�0�0�0�0�0�0 1(101<1d1p1�1�1�1�1�1�1�12 2H2h2p2x2�2�2�2�2�2�2�23(343X3d3�3�3�3�3�3�3�3$4,444<4H4p4x4�4�4�4�4�4�4�4�4505<5`5h5t5�5�5�5�5�5�5�5�5 6646@6d6p6�6�6�6�6�677787D7h7t7�7�7�7�7�7�7�7�7�7808<8`8l8�8�8�8�8�8�89949<9D9P9x9�9�9�9�9�9::::$:,:4:<:D:L:T:\:d:l:t:|:�:�:�:�:�:�:�:;; ;,;T;\;h;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<x<�<�<�<�<�<=4=@=H=h=p=x=�=�=�=�=�=�=�= >,>P>\>�>�>�>�>�>�>�>?$?0?T?`?�?�?�?�?�?�? p �  0 0D0P0t0�0�0�0�0�0�0�01<1D1L1T1\1l1x1�1�1�1�1�12,282\2h2�2�2�2�2�2�2 3333D3L3T3\3h3�3�3�3�3�3�34444<4H4p4x4�4�4�4�4�4�4�4�45585D5h5p5x5�5�5�5�5�566<6H6p6�6�6�6�6�6�6�6�6�67747@7d7l7t7�7�7�7�7�7888$8L8X8|8�8�8�8�8�8�8�8�8 9999 9(90989@9H9P9X9`9h9�9�9�9�9�9�9�9 :(:0:<:d:l:x:�:�:�:�:�:�:�:�:�:;;;;$;,;4;L;X;|;�;�;�;�;�;<<<<H<p<�<�<�<�<�<�<�<�<�<�<�<=0=8=\=p=�=�=�=�=�=�= >$>0>\>�>�>�>�>�>�>�>�>?(?0?8?D?l?x?�?�?�?�?�?�?   � �  0<0H0P0p0|0�0�0�0�0 1101<1`1l1�1�1�1�1�1�1�122@2H2T2|2�2�2�2�2�233<3H3l3x3�3�3�3�3�34,484\4h4�4�4�4�4�4�4 5@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�566<6H6l6x6�6�6�6�6�6�6�6�6�6 777$707\7|7�7�7�7�7�7�7�7�7�7�78$8,848<8L8T8\8h8�8�8�8�8�8�8 9949@9d9p9�9�9�9�9�9�9::<:\:d:l:t:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;@;L;p;x;�;�;�;�;�;�;�;<0<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�<==8=D=p=�=�=�=�=�=�=�=>><>D>L>X>�>�>�>�>�>�>�>�>,?P?\?d?�?�?�?�?�?�? � X  0 0D0P0t0�0�0�0�0�0�0�0�0$101T1\1h1�1�1�1�1�1�1 2,2T2t2|2�2�2�2�2�2�2�2�2 3 3@3L3p3�3�3�3�3404P4p4�4�4�4�4505P5p5�5�5�5�5�5606L6P6p6�6�6�6�6�6�6�6�677$7H7T7\7�7�7�7�7�7�7�7�7�7888X8d8p8�8�8�8�8�899(9H9h9�9�9�9�9:(:H:h:t:�:�:�:�:;; ;X;x;�;�;�;�;�;�;�;<8<X<x<�<�<�<�<�<=$=0=X=x=�=�=�=�=>8>T>X>x>�>�>�>�>?(?H?T?`?�?�?�?�?   � $   080X0x0�0�0�0�0�0(141@1d1p1 � x   `2h2`577 7(7,7074787<7@7D7H7L7X7\7`7d7h7l7p7t7h9�9�9�9�9�9�9�9�9�9�9�9�9::::$:,:4:<:D:L:T:\:d:l:t:|:�:|?   �   x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,202<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�243\3l3|3�3�3�3�3�3�3�344044484<4@4D4H4L4P4T4`4p4t4(5,5 <H<l<�<�<�<=(=D=d=�=�=>X>�>�>?4?\?�?�?�? � �    040h0�0�0�0�0181X1|1�1�1�12@2h2�2�2�23p3�3�3$4L4p4�4 5d5�5�5�5 6h6�6�6 7�7�7�78x8�8D9l9�9�9 :�:�:�: ;h;�;�;<�<�<=4=`=�=,>P>|>�>�>�>�>?4?X?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      