MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ��P�یP�یP�ی�2�Q�ی]��N�ی]�:��ی]�;���ی�m�S�یP�ڌ�ی�:�J�ی��Q�ی��Q�یRichP�ی                PE  L [ǵZ        � !    b     �.                               �         @                   `� [  � (                             ��  �O 8                           8 @              �                          .textbss                        �  �.text   x                        `.rdata  �Y  @  Z  "             @  @.data   �_   �  2   |             @  �.idata  �         �             @  @.reloc  l�     �   �             @  B                                                                                                                                                                                                                                                                                                        ������v ��� �l� �'� �� �� �. �� �` �> �� �f ��1 �X ��� �{ �V� ��o ��� �� ��I �ͮ �xr ���
 �>� 驒 �) ��� �z� ��	 �` �+l	 � �� ��� �gl �� 魋 �f ��� �5 �)� �d� ��]
 ��� �uG �0= �; �f� �1$ �< �7� ��
 ��� � �� �~G �	� �d�  �O� �� ��S �@_	 � ��I �& ��r	 � 钄 魁 ��� ��a
 �� �� �� ��� �� �%� �0� ��� �FF	 �� �l) �� � ��	 �� ��" 鎋 鉟 �� �?� �J  �e& �� �j ���	 ��� �L� �� �; �� �� �c� �� �Y �$� �ϡ ��  �J �� ��x �f �� �\! �w �j �� �h� �j �# �� �� �
 ��� �� �p� �˫ ��� �� �l} ��- �R� �� �� �� �^� �9� �.e ��  �Z� �uQ ��H �� �v� �� �< ��� ��5 �ͬ �hO �c� �^r
 陘	 �$� �_c �z�	 �5� �0� �k5 �C �q� �l$ �	 �r& �� �" � � �7 �� ���	 �
d �%D �P ��� �&� �1; �c �C �� �� �c �#� ���
 �Y �T �o`	 �:C �e� ���  �z �� �c ���
 �� �r� �m� �- �S� �>@ �# � �//
 �N �5� �Xd 黇 �F�  ��O
 �| 
 �c �2� �� �xj �n �~� �� �� �� �j �%� �p �+d
 �6� �1�	 �l� �� �r� �-< �x� �33 �M �� �4& �O� �:� �u� ��	 �k- �' �1�
 �L� �7Q �b �]�
 �(6 � �c �)� � �� 骸 �U� �� ��Q �&� �qi �O ��� ��a �q �S �Q �. �	 ��� �o� ��  �5� �@� �� ��  �qM �<U �Ga � ��" �8 ��
 ��� 鹡 ��� �O�	 �
X �%$ �p�  �[$ �� �� �̥ �' �� ��o �H� �3a �^B �n �$� 韛 �Z �5�  �� �� �&� �] �LY ��o 邽  ��� ��� �S,
 �� ��� �
 ��Y ��\ �u�	 � � �� ��� �y � 駯 �� �- �h� ���	 �n� �iP �� �C
 ��	 �U_ � � �{� �V/ �qp �] �W� �L �=� ��` �A
 �nm �9� �4� ��Y	 �� �� �� �� �� �U| �\4 �R �RI 魢 �` �#� � �� �D �O� �*U ��S �0 �[	 �V� �1� ��b �a �b� �% �" �# �� �Yv �f �� �ڨ �c ��| ���	 �6� �qi ��  �'�
 �RM �m% ��� �s� ��
 �" �� 鿍 �
� ��� �] �[\ 閧 ��j
 ��B ��2 �bI �� �Ȧ �C� ��� ��t 鄤 �O �ʤ �uJ ��� �{�	 �$_ ��� �<� ��A �r� �� �� ��i �~� �9	 �d� �� �ڲ �E  逜 �{ ��  �!� �:	 �g�  �B 魇 �x_ ���  ��7 ��� ��� �ߪ 銰 �Et ��3	 �S
 �vU �C �, �g? ��t �M �x ��  ��J �i` �h �?g �e �� �0u ���  � �q4 �_ ��^ �R�	 �}� �� �3� �n� �� �D1 �O# �:L ��c ��a �[� �= �a�
 �<� �S �2� �=C ��� ��2	 �Ni �	�  �4V �?8 �:( ��0 �p� 鋴 � �� �w 问	 �B< ��� �ؒ �N �&^ � �� ��e
 �� �E� ��  �� �&8 �q� ��K
 ��5 �Y ��k �� �# 鮓 ��p 锗 � �5@ ��W	 �0� ��� �v� �q> ��� ��� �z �}� �8� �d �N� � ��� �� �ڴ �M\ �P� ��� �&b �q� 鬺 �gX	 �' � �X1 �s�
 �� �9} �Ĭ �]
 � ��K ��\ �{� �? 顽 �| ���  颸	 �=�  �8� �C� ��� �y@ �D! ��? �j� �� ��? � �vH
 ���  �/ ��	 �2� �]� �� �# �n� � ��z �_ �j9 �� 逬 �ۓ
 �E
 �19 錤 � �+ �M� �H 飐 �>� �y �; ��� ���
 �e� �pZ ��/ � �Ѭ �,* ��� ��% �7 ��� �� �nk �YF �T� �/> �:� � � D
 雝 醖 �!� ��Z ��# ���  �M� �Ȇ ��P �N� �� �TN �O �� �Ձ �� ��V	 � 
 �A4 ��� �7} �J �}� ��� �F �>� �9 �$3 �/9 ��� � ��^ ��H �&� �[ �: �� �2 �( �h� �oZ �>� �٢ �$) �/j �zG �� �. ��E ��x � 鬥 � �� �]u �8 �� �� ��: �Դ	 �� ��R �E�  � � �k� �f
 �1� ��J �w�
 �� �m0 �� �c
 �� ��� 锢 ��� �
�	 �� �� �+�  ��� �� �� ��j ��� 齏 ��N �� �N0 �iG �t� ��� �Z� �2 ��� � ��: �� �l� �I	 �� 魕 ��  ��_ ��� �i= �O 韸  �Z� ��� �P� �{�
 �j �
 �|� 鷎 �� �^ �� �� �
 �9� � �/ 骷 �8 �0
 �ˬ
 �� �Q�  ��� �G� 钮 ��	 �x=	 �sY �h �g ��
 ���  ��� �5� ��L �k� ��	 �+ �,� �� ��� �� ���	 �� �~� � �$z �n �T	 ��� �p ���
 閌	 � �/ �'� �� ��� �| �gX �^� �9�  ��C
 ��  ��� � � � �{  ��� �O �L �Ǯ �hX �- �, ��� �Y �  �� �ϩ ���  �e� ��] ��b
 �� �a- �� �w< � �� ���  �3� �� �� �$E
 �� �� �� �@f �r ��W �q�
 �<@
 �צ �҅ ��	 �h� �s� �� �� �t �/� 銂 �� ��P ��	 �W �^
 �L� �� �RV �E �
 �� ��� �R	 �t� �_E �* �%�
 �pI ��� �4 �� ��6 �W
 �B1 �]� �; ��+ �P	 驯 鴬 �� �Z� � �W �;w �� 遍 �L3 �7 ���	 齾 �� �q �n�
 �� �d' �� ��  �� �@�
 �u �V� �B	 �l8 ��	 ��  ��K
 �� � �P	 �ɀ ��, �� 銏 �� �� �{�	 �f �1� �� �'� �� �--
 �Ȉ 郻 ��� ��k	 �D� �o�  �ڍ �5]
 �p�  � �	 �� ��� �T �rE �}{ ��	 �C� ��� ��� �� �O/ �� �ŕ 鰁 �[ 鶯 �!� �� �׆ ��� �� �x�  �#� �. �9 �$� �/^ �u �5�
 造	 �� �fC �� �� ��2 ��� �-7 � �C� �� �� 锪 ��F �j �E� �� �˥ �	 ��� �� �G�  �b�
 ���  �x` �c �n� ��� �t} ��� �Z� �5 ��Y �� ��[
 � ��� �wk �Rh	 鍼 �� � �N�  �IL �� ��� 隷 �uD �0 �
 �� ��r �|+ �W �& 鍹 ��	 �� �� �&	 ���	 �_� ��� �� �@}	 ��6 �� �!�
 ���	 ��	 �� 鍙 �� �ӽ �^�	 ��
 � �O| �# � �p� �� ��� �1� ��, ���
 �� ��  ��+ ��O �� �)� �t# �O� �Z� �U� 鐰 � �6� �Q �\� �g� �4 ��# �H �S
 �� �i� 餠 �_2 �j	 ��! �н �� � �!� �l� ��l �b� �}� �H� �� �n� �� � �� �*� �� �@ �k� �� �� �l* 闩 �� � �x8 ��  ��	 �p� �d� �/H �j �E� �`�  �+�
 �V �!� �| �Ƿ	 �| �]; �� �# �nE �yy �d
 �?m �� �e� ��3 �k� �vN �Q� �̲ �L � �=� �X 鳎 �n� �� ��{ �W �j� �5� ��k �{5 � ��C �,S �w� �b ��. �hq �- ��H �� �- ���
 �
@ �5 頫  �<
 �� �B �,{ ���  ��  �-� �, �S� � ��� ��x �O} �j�  �� ��s �;. �� �1; ��� �7� �b �]� �hh	 �3y �5 �٤ �$; �? �:t �u) ��Q
 �K� � �qx �� �� ���  �݃ �(F 铥 ��H	 �	�  ��a �o�  �*� ��� ��  �� �� ��� � �  ��	 ��� �(p �C �n �� ��S ��I �� �U
 � P	 �m �f� �AM �L �H 邟 ���
 ��� �� � �� �t[ ���	 �� � 鰃 �P �� �A ��  �w
 �<� ��| �ظ
 �
 �� �� �( � �Z �� �p�  �� �H �| ��  ��� ��� �. �g �3? �>� � �$� �O� �
� �� �� ��B �b �!H	 �| ��� 顭 �]� ��6 �� �S
 �i�
 锑 鏄 �j�  �e� � � �+f �v
 ��C �� ��g �� �-� �� �% �N� �o �t, �: �z �E  ��N �
 �� �| �T
 � 邴 ���
 ��M 飃 � �yN
 �� �Om �*
 ��
 �0� �F	 �) �q� �\� �g  �R? �� �� �r �w �� ��? �� ��  �� �`�
 �+� �� �KN �l� 闔 钝 �=�  �(A �#� �n7 �� ��` ��  ��M ��	 �0X ���  �6�
 �� �� �� �b� �� �(� �� �n� � ��� 韾	 �z� �e�  � �;� �v> �� �|� �Wq 鲂 �}� �HG	 �- �^q �)� 鴁 �O�	 �*8 ��K � ] �{W �F� ��  �l� �h ��3 �� ��  ��	 �n� 陵 �d� �h �Q �E �Щ �K0 �� ��� ��f �6 �� ��  �� �� �� ��	 �)	 �� ��d �z ��� �;2 �։ �As �� ��0 �2� �}� �dK � �� �	� �D�	 �o� �:� � �@ ��� �F ���  ��� 闙 �� �� �h �#� �� �٫ ���  �O< �n �9 �� �;� �Q
 �q� �< �. �J �-� 騪 �U �N�  �
 �d� �� ��� �| �P*	 �+� ��- �q�	 ��� �+	 �"� �4 ��� �iJ ��w �� 餘 ��� �� �0 �0� �[; �� � � �}
 �rx ��� �( �3& �n� �)� ��I �s ��  �� �S
 �� �V �g �� �'N �� �� �F �cJ �a �	� 鄆 鿝 �"
 �� �  �+� ��� �� �|� �� 鲋 �I �X�
 �H �ށ �)� �4
 �� �ʺ
 �� �  �| �� ��G ��  �p �r  �-~ � ��H 鞅 �i~ �� �n ���  � �P�  �ۥ	 �6 ��� �̧ ��
 ��Y �  ��N �� �^�
 ���	 �D� �� �5 �Es �0� �\ �f ��{ �� �'� �2� �-� � �s�
 �N�
 �4
 ���
 鿩 �� ��� �@� �� �} �� ��� �׾ �� ��
 ��Z �C�  �>�  ��  �� 鏆 �j� �� �`� �� �6� ��
 �\� ��C �� �}'	 �(� �z �� �� �t �Ot ��� �? �`� �+�
 �� �!� �� �g�
 �� ��t ��M �s| �N ��� �I �/�	 ��� �� ��� ��H �  �� �\}	 �� �B �}� ��� 鳾
 ��
 �h ��	 �" �B	 �+ ��F �[� �<
 鑣	 �,� ��  �b ��E 騤  ��	 ��  �Y �TE �, �
� �ej �@� �;� ��� ��  �L� ��n �2�
 �=& �� �s0
 �>� ��\ �4
 �o�  �| �5 ��3 �+� �f � ���  �� ��  �=� �X� �q �5 �� �� �	 �ZJ
 ��� �� �OF �� � �B �g+ �2q �� �x�
 �C 龥 �T �� ���
 ��A
 ��� �v �< �6L �1� �M ��� 鲙 �� �� �S�  ��� �� 鴾 �V ��� ���  ���  ��# �&�  �a� �} ��, �� ��  ��� ��� �f �	� �� ��v �ڱ �q ��U �sF �3 � �K �7� � �=� �x� ��	 �~  �Y� �$� 韫 �*` �u< ��, �x �6W �Ѱ �� �Ǧ �R� �� �8m	 �� �� �y, �bE ��� �J{ �Ű ��( 雛	 ��� �Q �� �W� �� 魺 �� �	 ��. �Yt �� �_� �J �� � � �+� �Fx �1} ��- �G �2� �� ��W �l' �^  �9� �� �O� 麮 ��� �p� ��� ��' 遻
 �� �W�  ��5 �=	 �� ��<	 鮠 ��o �� �o� ���
 �} �0�  �KS �&�  鑺 � � ��A	 �� �X, �� ��� � �9
 �� �J� �5� �	 ��  �� �� �l= �k �2� �ݕ 阋 �� �N �	 �a �� �::
 �U ��  �k� 鶲 �� 錦 �� ��� �2 �� �# �� � �q � �z� �5� �p�	 �K  �&G �Q� ��
 �# �2�	 ��� �\B �#�	 �~' �9�  �T� �� �
3 �3 ��4 �� � ��  ��� �d �� �� �H� �S�  �~� �ّ �D~	 �� ��� 饑 �� �� �F�	 �Q� �L� �j �P� ��� �x� �#� ��r ��� �� �/� �
? ��C �� 髇 馌 ��� �~ �'� �b� �Mp	 �� �S� �.� �) �� �?� �j ��� � >	 �5 �&� �q� �\� �w� �2� �m= ��% �3� �� ��� �B �� ��� �E� �0� ���
 �V ��  �$ �. �� �Ͱ ���  �3� �>4 ���	 �T� �_� � ��  � � �;� �& �Q ��� �W �r�  �� �z �� 鮢 �y� �H
 �_ � ��  �p
 � ��H �An �,� �N �3 ��" �( �C! �� �	� 鴌 韱 �f �E� ��� ��k ��  �Q~ �� �{@ �ra �-+ 鈟 �� �>� 鹩 �T �o� �J� �5� �� �� �fH ��2 �|} �g� ��� �}s �8 ��Y �~K �i{ �$� �?� �� �e1 頴 ��� �� ��~ �\g ���  ��� �] � �c� ��H �� ���	 ��� �
� �� � �ks �V�  �� �� �GG
 �� �M4 �8 �SP �^�  �y� �� �o		 �j� �ul �� �k,
 �֊ 鑁 �;	 �7J �҆ �M� 鸄 �@ ���	 �p ���  �� � ��� �0�
 �k�  ��� ��	 �1 �� ��� �%@ �H� �ã  �^ ���
 锺 ��{ �J� �%� � � �! �O �� �� �Wo ��� 齈 ��� �� �^j �iD �Tu ��� ���	 �E�  � �  ��� �fC	 �� �' ��` �Rb �> �� �3� �> 驆 �dq 鯰  � ��� �2 �KM �v� �A� ��P �7 �� �}�  �X� �C�  �� �I; ���  �� �& �� �� �Kb �� ��  ��� �g#
 ��  �" ��
 �� �no �� � �h ��� 鵹 ��� �g �� �A� ��  �7� � �-� �� �:	 �n� �)A 锐 ��� �z ��# ��
 �{ �� �A�  �l  ��I ��w �� �s �C# �� 鹼 �f	 �� 銌 �U< �C
 �e �ֱ �!�  ��< �g� �B
 ��D
 ��W �s$ �� �i* �D� �e 麊 �%� �r �3� �;	 ��
 ��
 �' ��� �� ��� ��u 鎋	 ��� ��� �� ��m �� ��� ���
 �& �� �� 釕 ��
 �-Y	 �� �z �^
 �	Z �$� ��) �*B
 �E2 �r �۹	 �� �q[ �|? �) �� �m �H` ��
 �^� �� �K ��  �ڤ �Y � h 鋘 ���  �< �� � � �� �	 �]	 �~o ��: �z �� ��� ��C �`4 �� � ��> �l�
 ��
 �r� �]� �� �c �~ �O 鄎 �߱ �� ��  �� ��k �F  鱲
 �\� �g� �� 鍒  ��� �� �>k �in � �� ��)	 �u� �	 �+� �N ��  �Z �ǜ �% �-�
 ��� �< ��
 鉂 �t� �} �*n �%j � �� �: �e ��  �w� �R �� �H\ �c� �^� � �t� �� �Z� �5W ��] �: �&�	 �!� �� 鷳 �g 鍧 �(� �#� �� �� �� �� ��
 镄 �@ ��� ��) ��O �L�
 �� �� �=& �D �d �6 ��	 �� �� �� �e�	 �0  铘 �� 鱕 錧  �G� �R�	 �� ��{ �~	 �~� �& �d� �O�	 障  �� �� �K� �f� �0 �� �H � �m �� ��� �Nx �)	 �T�
 ��| �:� �%�  �@�
 �+� �� �A� ���  �G�  �J �mb �Xn ��  �n� 鉊 �Է ��� ��� ��V �0�  ��  � ���
 ���	 �7�
 ��[ �m� �h* �c/ �~ ��3
 ���  �� �C �5:	 �0� �{� �v� �! �� ��@
 �B� �7 ��4 �s� ��7 �u 餾
 �9 �J� � ��J
 ��
 �&� ��� �<' �� �Bk �� ��0 �3 �N� �i �� �o'	 �:� �� ��a ��	 �F� ��� �\ ��  �_ �]& �� ��� �>� �3 ��6
 鯮 ��� �u� �� �kY �J� �qk ��� �g� �& �� 阦 �� 鞸 ��
 ��� ��,
 �j� �E�	 �p�
 � ��j �1� �� ��� ��� �6 ��U ��	 �� �Ɇ �[	 �?�	 �J	 �� �{ �۵  ��
 �Q] �y �7� �F �-4 �� �#� �~p �)�
 餜 鏧 �j! �u� 逴 ��z �6 �a& �, ��� �G �-� 鸋 �� 鎚  鉳 �4 韉 �J� ��
 �P� �[J ��� �A �l� ���  �«
 ���	 �X� ��  鮞 �9� ��� ��{ �
� �} �� �� ��  �� ��g �� �2�  �=� �(� �S� �> �z �d� �?� �J. �U� �P� 鋹	 �V� ��0 霤 ��� �� �{ ��6 �s� �% �)� �D? ��	 �� 酐 ��� �� �f] �Q! �|
 ��
 �� �� ��� 鳤 �~� �Y� ��� �OY ��� �z	 �� 黚 �fj �� �,. �W� �� �m �ȁ �� �� �G �$�
 ��e 銌 �� � � �� �v� �� �l �e ��` �m� �4 ��
 � ��� �$� �� �z� �o ��� �+� �1 �� �� �� �R� �}�
 �m � ���
 ��� �t� �q �.4 ��] �Р �+K �� 顒 �,	 釣  �B? ��	 �x� �� �.� �i� ��3 ��" 麄	 �E �� �� �� � �w 駑 �\ �-� ��  �Ӹ	 �>� �� ��� �o!
 �JJ �e' � d ���	 ���  �� ��	 �w[ �� �) ��� �b �^�  �YO �d� � �j �3 �P% �� �� ��* 霴 �gI �� �]T ��	 �֑ �ޯ �c �$� �O� ��� �� ��  ��� �+ 韑 ��` �Wc � � �h� �� �~ ��� �4a ��
 �� ��
 ��, �k� �F� ���  �\� �� �r� �m� � 郠  �n� ��	 ��� �" �
 ��
 � � �2 �& ��
 �\�
 �� �2 ��D	 ��U �#p �n �9�	 �dw	 �\ �
 镣 �@g ��� ��� �Q� �� ��� �R� �� �X�
 �S& ��k �y� ��+ �� �� �N ���  �{� ��� ��c �<_ �7� �҂ �# 鸎	 ��f �*� �I� �� �` �� �e7
 �p� 雺 �z �P �\� ���
 � �=� �0 �� �.� �I �D� �� ��� ��� �0-	 �K� �V �� ��4 �w ��  �\ �8K �s �� �9�	 ��
 �o� �
� � � u �;� �v� �A� �|� ��  �@ �M
 ��� �� �~D ��  �D! ��� �j� �U� ��% �[P �� �" �l� �� �2� �]( �hg �� �~ �i �� �" �Jt �2
 �p� � �o �� 霩 �g ��	 �M� �h�	 ��V �q 鹿 ��! �| �j� �%4 � � �� �&	 �� �L+ �~ �2 �ͽ �H� ��� �� 鉮 �4�  ��� �z�	 �� ���  ��
 �&E �" ��� �7( 钑 �Z �ȸ �#% �� �Ig �� �2 �
� � 頓 �;� 馄 �� ��	 �7� �" 靤 �� ��� ��
 �V �t�  �ڽ	 ��O �� �x ��P �6�	 � ��	 �7� 钴 �-� ���
 �� ��� �� �* �� �� �� � �k�
 �6S � �t �� �r� �� �(� �p �~S �Y�  �d� �/� �� ��6 �0� �K9	 ��(
 �! ��Z 駅 颼 � ��w �c�	 ��  �y� �� �	 �Z� ��# �  �[� �M �P�	 �|� �i �"�	 �� ��+ �c� ��� �� � �o� � �� �0�  �1 �v� �1� 錿  �Ǥ � �̀ �o 鳆  鞯	 � ��� �o~ �*� �
 � d �� �@ ��� �,� �, �"�	 魾 ��� �#� � � �� �_� ��� ��> �8 �{)
 �6)
 � �+ ��  �R
 �=� �Hv �#P �>� ��b ��^ �ϖ 麭	 �u| �� �Z �o	 �Q$ �̠ �Wm	 �"� �m �8� �3� � �) 鴣 �_� � �5' �% �+ �6� �	 �܇	 �7�  �2� �	 �� � �n� �)� ��< ��a �h �+ �>+ �[� �v ��� �<| �x ��q �� �h� �c� � �S	 �� �� �( �} � [ 雏 閞 �1 �� �W� �� 靑 �� ��j ��  �iu �� �O� �Z�
 ��� �p� �� �v� �!� �<� �g� �" 鍴 ��� �#� �n+ �I! �� ��� �z�  �Ew �- �;� 醧 �� �ܪ �W[ ��� ��&
 �x� �1 鮦  �I� ��B � �j� ��V �@� �"� �6O � �&
 �'� �;� �'� �� �� �n� 鹹 �� ��� �� �� �[ �˯ ��+ 鱍 �� �Ǖ �r� �]� 鸶 �ì ��O �Y> �tQ	 �� ��` 镄 �P�  �S �V
 �# �
 �7� �r� �M> �q �d �� �)� �4M �} �ZY � �V �_� 醮 �i ��� �<� � �O �P	 郑 鎑
 ��z ��k	 �O� 隀 �� �ݵ ��  �* �Ae �|� ��6 �2�  �=�  �� �� �} �Y� �D� �OY ��
 ���	 �pK �� 
 ��B �=) ��	 �� ��
 �M �� �Cv	 �^h �ٷ �dw �p
 �*� � ��� �+ ���	 �Q �|�	 ��	 �r= �ݿ �H � �ޠ �Y� ���
 �� ��z �� � �7) ��� �� �O 駥 �" ��  �H1
 鳂	 �~ �9� �T� �y �J� �� �px �;� ��0 � �lN ��Q ��` �m� ��� 鳖 �N[ �iq �tK �v ��
 ��� �� ��&
 �v
 �q� �� �g �� �]� �X� ��� �~� �	� �D� �/� �*K 鵔  頺 �b �6� � ��� �  颕 �=� �8u	 �� ��b ��  �� ��� ��� ��  �p� � ��� 鑾 �� � �R: 齃 ��L �s�	 �l ��� �x �?N �
 ��% �`4
 ��� ��w �� ��" �g� �t �=�  �� ��� �e �I� �$ ��� �z] �UB 逞 �� ��	 額 錷 �� �& �B �x� �� �� �9� �D!
 �� �g 饿 �pE �;� �W �1� �z ��	 �� �=� ��v �� � �)!
 �T� �_� ��" �U� �l �KZ �� ��	 �\� �� �� �{ �"
 ��  ��� ��V �D� �o� �*D �uC �PB �u
 �w �� �� �V ��C	 �-W ��  �#� �� �)� �� �� �H% �u� �p� ��  ��� �Q� �] �� �b� ��x ��M	 �æ ��D �ɯ �Tf �5 �
� �eM �@} �� �&w	 �Q� �� ��� �b% ���  �h� ��� �Ns ��L	 �� �o�  �% ��� �0� ��	 �� ��� �<{ ��? �� �]� 鸿 �Z �N� ���  �4�  �O� 銫 �E� �$ ��q	 �& �1J �L ��m �2� ��� ��$ �� � �y� ��� �� �*� �u�  �� �۠ �& � �l� �# ��� �r ��%
 �ó ��� �� �/� �� ��  �� ��R �k	 �F� ��� ��J �G� ��� �-� �y �S�  �>�  �y� �$ �8 �jg �
? �p� �k` �f� �] �,� �&
 �� �]  �x� �
 ��� �9� �Է �o	 �� �] �0a �� �d �� ��) �G� �r �r �� �s� �N
 �Y�	 ��� �� �j� �E| �@� �K� �L ��� �L �� �R �o �� �S� ��� �i� �� �x �J �eU
 ��� �;M �6� ��* �L 闺 �� �-� �m	 � �~" �T �d�	 韹	 �J� 酏 �p�  �ۤ �V� �12 �� �G�
 �� ���	 �(\ ��� �d �ɠ ��	 �?� ��� �� �P� �K �� �A
 ��s �� �� �m� �X�	 �3V �~� �i�  �� �N ��s	 饏 �! ��| �� �_ ��� ��a ��	 ��) ���
 �Ø �Nk �9� �ė ��T ��� ��	 �P� �� �	 �A�	 ��n �� �R�	 ��h �(� �! ��Y ��I 餧 �O6 �:� ��� �0� �Kd	 �f� ��� �,K ��� �! �}� �آ �C/ �nx  �v ��M ��E �
� �� � ? �� �f� � �,C �Wk �b� 齆 鸣 �S^ �~� �	q �6 ��� ���  ��	 �� �\ �� �A� 霕 �'� ���	 �]� �X� �S( �.�	 �H �$1 ��� �0 �5� �0 �T�	 閫 �� �\) �'n � 鍓 � ��}  鎩  �� �$i ��> �� �e� ��
 �{� �F� �љ ��	 �W� �� �� �S �S� �~�  �-
 �� �?I 骮 ��  �@F �{� �&/	 �q� �\ ��! �b� �* ��� �S� �� �)� �D� � �jj �� �� �˫ �vk � �|� �G� ��n ���
 �(�	 �C� �% 陓 �t
 �?� 骉 �E ��J �[& �	 ��� �\n 闡	 �� ��� �H� �� �n	 �P �tN ���
 隝 �#�	 �	 ���  �� � �<$
 问 �1 �� � �� �N� �� �D� �O� �zj �� �`q ��� �&p �!} ��T �g#
 �� 鍰 �(� 铒 ��% �y� �8 �_# �� ���  �p� �� � �� �\� �4 �%
 �}$ �� �	 �n�  ��F � ��� �*� �� ��� ��s �fs �o �,U �
 �% �=p ��%
 �� ��o ��� �� 韚 �: 饶 ��  ��� � �!� �i �V �� � ��n 鳓 ��b ���  �ԙ �� ��� ��� �� �{	 �L ��z �̇ ���  ��� ��� �x� �|  �.� �	o �$� ��� �j� ��$	 � � �� �&� �1� �\S �G�  �� ��� � ��� �^  �� �� �� ��D �o �Pd � �d �!� �F 駰 �b� �� �H1 ��� �~B 鉏 鄬 �Ϭ
 �z�
 ��� 鐚 �+t ��� �1�  �,� �� � �m� �8L 飛 鮭 鉯
 �D.
 ��� ��
 �e� �� �K� �Ɲ ��	 ���  �� �R� �� �� � �n� �9 �ď �O 麌 �5� � � �, ��  ��| �e �7 ��	 ���  �� �c* �  �� �t� �ϱ ��/ �� 鐊 �� �V� ��	 ��X �� �b| �R ��� � �ι �yz �Դ �/� �ڦ �Ŏ � � � �&� �A�  �� �- �r  �=� ��� ��� �~Z ��� ���
 �o� ��  钩	 �`p ��� �v} �� �� �} �Ҍ	 ��t �� �C
 �� � �4� 鏶 �J� �U� �  �� 馚 �Q� ��v �u �� ��2 �8� �3� �> 驛 鴽 �g �J� �� �`% ��? 香  �� ���	 �'� �2 ��
 ��J �c �n� �� �dz  ��� ��  � � � �Y �K � �9 �5 �r� ��� �Ȝ �3O �^  ��H ��� � �v �� �@� �
 � ���  �l ��� �r� �}m ��D �ӓ �^� ��j �T�  �o� �e ��* �@� �;i � ��I 鬁 �W� �bt ��� �H� �& �n� ��: ��� ��: �:� �� �`< �[�  �v� �Q; �<j �g� �; �ݽ �(� 鳂
 �~� �	� �T� 鿩 ��� �4 �Д �;� ��� �1� �u 釃 �� �� �Hj �� �n �? �$ �OO �
� �k � �{� �f= �� ��  ��  �x �� � �#� �q 陜 �� �d �
� 镘 � 3 ��	 閝 鱢 �l� ��# 钽 �� ��  �sF �~k �ym �$� �� �: �ş �@� �+�	 醰 ��� �� �G� �r�  �-
 鈿  �C� �~� ��9 ��G �� ��� ��E �� �k �&
 ��� �LN �Ǽ  �� �E �� �s �.� ��� �� ��  �� �Ej �P� �;O �&	 ��� �l� �ף �j �Q �` �� �nV �I �4� �� � �� ��R ��^ � ��  �� ��_ ��L �}� 鸐 �c� ��	 �i
 �W �?d �z� �
 �Ђ �ۓ	 �~ �
 ��� ��  �� �=� �� ���	 �.� 鹦 �t �o� �jC �� �2 �k� �fu � �ܦ �h	 � ��
 �H� ��� �j �y 鴄 �
 �8 �E� ���	 �KJ �f� �Ѳ ��a �s �� �Mt 阎 �Û �� �Ij �� �/4 �:� �u�	 ��	 �M ��� ��� �<� 闗	 �R� �}� �J	 ��p �.�	 �	�	 �g 鿪 �z�	 饌
 �0{  ��� 馲 ���
 �|� �Ǒ ��� ��E � �8 �nL �9
 ��t �� �J� �e ��
 �� � �1	 �ܔ �G� �� �� ��j	 �� �>H ��� �_ �� �z �%	
 �p  髰 �l �� 騣	 �gI �k/ �=M �8� 飦 �~= �% ��. ���  �a �� � K ��b 馪 ��� �\I �v �C� ��1 ��P �2 �.� �	� ��K �� �*^ �P ��� ��  ��� 遺 �l�  � ��3 ��N �ȗ	 �3� �.� �� 鴶 �� �x �5� ���  �k� �vO �q= �� ��� ��� �� ��� 鳞	 �~� �YK 鄸 韖	 �f 鵸 �E �˜ �q� 顝 ��
 �w� �� �ͽ  �H_ �� �N� �� �� �ߩ �L ��� 項 鋄 �� ��  �� � ��> �=� 阄 鳶 �  �	 �dO �� �� �5� ��� ��� 馩 �a�
 �|P �� ��� �� �8� ��} 鮈  �	� �t� �_� �I 鵭 �� �;� �F �AB � ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   ���������ko��hP'�A�����_^[���   ;��j�����]������������������������U����   SVW��@����0   ���������Y��h�'������_^[���   ;��
�����]������������������������U����   SVW��@����0   ���������z��h�'�����_^[���   ;�誓����]������������������������U����   SVW��@����0   ������j ����U��_^[���   ;��U�����]�������������������U����   SVW��@����0   ������j ����:U��_^[���   ;�������]�������������������U����   SVW��@����0   ������j �����T��_^[���   ;�赒����]�������������������U����   SVW��@����0   ������j ����T��_^[���   ;��e�����]�������������������U����   SVW��@����0   ������j ����JT��_^[���   ;�������]�������������������U����   SVW��4����3   ������3���;���_^[��]��������������������U����   SVW��4����3   ������3���;���_^[��]��������������������U����   SVW��@����0   ����������S��h@(�}����_^[���   ;��:�����]������������������������U����   SVW��@����0   ������j ���膂��_^[���   ;�������]�������������������U�����g���h�(�||����]���������������������U�����vk��h�(�L|����]���������������������U������U��h�(�|����]���������������������U�����yv��h�(��{����]���������������������U��j ����%R��]����������������U��j �p��R��]����������������U��j �����Q��]����������������U��j �t���Q��]����������������U��Q3��E���]����U��Q3��E���]����U��m��}��]������������������U��Q3��E���]����U�����j��h)��z����]���������������������U�����~T��h0)�z����]���������������������U�����u��hP)�z����]���������������������U��j �����P��]����������������U��j ����P��]����������������U��j ����P��]����������������U��j ����eP��]����������������U��j ����EP��]����������������U��j ����%P��]����������������U��j �p��P��]����������������U��j �����O��]����������������U��j �t���O��]����������������U��hp)�Fy����]���������������U��Q3��E���]����U��j ����zh��h�)�
y����]�������������������U��Q3��E���]����U��Q3��E���]����U��Q3��E���]����U������g��h�)�x����]���������������������U�����>R��h�)�|x����]���������������������U������r��h�)�Lx����]���������������������U��Q3��E���]����U��Q3��E���]����U�����&g��h*��w����]���������������������U�����Q��h0*��w����]���������������������U�����)r��hP*�w����]���������������������U��Q3��E���]����U��Q3��E���]����U�����vf��hp*�Lw����]���������������������U������P��h�*�w����]���������������������U�����yq��h�*��v����]���������������������U��Q3��E���]����U��Q3��E���]����U��Q3��E���]����U�����e��h�*�v����]���������������������U�����P��h�*�\v����]���������������������U�����p��h+�,v����]���������������������U��Q3��E���]����U��h0+��u����]���������������U��D��{��hP+��u����]���������������������U��Q3��E���]����U�����d��hp+�u����]���������������������U�����O��h�+�\u����]���������������������U�����o��h�+�,u����]���������������������U��j ����eK��]����������������U��j �\��EK��]����������������U��j �`��%K��]����������������U��j ����K��]����������������U��Q3��E���]����U��Q3��E���]����U�����c��h�+�\t����]���������������������U������M��h�+�,t����]���������������������U�����n��h,��s����]���������������������U��j ����5J��]����������������U��j ����J��]����������������U��j �����I��]����������������U��j �����I��]����������������U��j ����I��]����������������U��j ����I��]����������������U��j ����uI��]����������������U��j ����UI��]����������������U��j ����5I��]����������������U��j ����I��]����������������U��j �����H��]����������������U��j �����H��]����������������U��j ����H��]����������������U��j �x��H��]����������������U��j ����uH��]����������������U��j ����UH��]����������������U��j �p��5H��]����������������U��j �|��H��]����������������U��j �����G��]����������������U��j �����G��]����������������U��j �t��G��]����������������U��j ����G��]����������������U��j ����uG��]����������������U��j ����UG��]����������������U��j �t��5G��]����������������U��Q3��E���]����U��Q3��E���]����U�����_��h0,�p����]���������������������U�����J��hP,�\p����]���������������������U�����j��hp,�,p����]���������������������U��j �0��eF��]����������������U��j �4��EF��]����������������U��j �8��%F��]����������������U��j �<��F��]����������������U��j �D���E��]����������������U��j �@���E��]����������������U��j ����E��]����������������U��j �p��E��]����������������U��j ����eE��]����������������U��j �t��EE��]����������������U��j �H��%E��]����������������U��j �L��E��]����������������U��Q3��E���]����U��Q3��E���]����U�����]��h�,�\n����]���������������������U������G��h�,�,n����]���������������������U�����h��h�,��m����]���������������������U��j ����5D��]����������������U��j �p��D��]����������������U��j �����C��]����������������U��j �t���C��]����������������U��Q3��E���]����U��Q3��E���]����U����   SVW��@����0   ������E���Ex��M�U;��G����EE�E��_^[���   ;��,�����]� �����������������������U����   SVW��@����0   ������_^[��]������������U����   SVW��<����1   ������E��<�����<���t�����^C����u3��3�_^[���   ;�艀����]�����������������������U����   SVW��@����0   �������&�����u3���   _^[���   ;��/�����]�����������������������������U����   SVW��@����0   ������E;Et��EPj �MQ�Zl����_^[���   ;�������]�����������������������������������U����   SVW��4����3   �������E�    �} u� �}�w�EP��Y�����E��}� u�TP���E�_^[���   ;��?����]�����������������������������U����   SVW��4����3   �������E�    �} u�&�}���w�E��P�XY�����E��}� u��O���E�_^[���   ;��~����]���������������������������������������U����   SVW��4����3   �������E�    �} u�$�}UUUwkE0P��X�����E��}� u�@O���E�_^[���   ;��+~����]�����������������������������������������U����   SVW��@����0   ������} t#��j �E��M���;���}���EP�L�����_^[���   ;��}����]��������������������������������������U����   SVW��@����0   ������} t#��j �E��M���;��D}���EP�̇����_^[���   ;��(}����]��������������������������������������U����   SVW��@����0   ������} tj �M�F?���EP�Y�����_^[���   ;��|����]�����������������������������������U����   SVW��@����0   ������} u�EP�MQhH]�e����_^[���   ;��F|����]��������������������U����   SVW��@����0   ������} u�EP�MQhH]�3e����_^[���   ;���{����]��������������������U����   SVW��@����0   ������} u�EP�MQhH]��d����_^[���   ;��{����]��������������������U����   SVW��@����0   ������} u�EP�MQhH]�sd����_^[���   ;��&{����]��������������������U����   SVW��@����0   ������E;EtE�EP�MQ�UR��}�����EP�MQ�UR�}�����E;Es�EP�MQh�]��c����_^[���   ;��z����]����������������������������������U����   SVW��@����0   ������E;EtE�EP�MQ�UR脍�����EP�MQ�UR�p������E;Es�EP�MQh�]�Ac����_^[���   ;���y����]����������������������������������U����   SVW��@����0   ������E;EtE�EP�MQ�UR�|Y�����EP�MQ�UR�hY�����E;Es�EP�MQh�]�b����_^[���   ;��Ty����]����������������������������������U����   SVW��4����3   ������EP��;���Q�p�������P�MQ�UR�EP�MQ�~G����_^[���   ;���x����]������������������������������U����   SVW��4����3   ������EP��;���Q�f�������P�MQ�UR�EP�MQ������_^[���   ;��Px����]������������������������������U����   SVW��4����3   ������EP��;���Q��Q�������P�MQ�UR�EP�MQ�U����_^[���   ;���w����]������������������������������U����   SVW��4����3   ������EP�MQ�h������;�����;���R�EP�MQ�UR�Nm����_^[���   ;��Ow����]�����������������������������U����   SVW��@����0   �������	�E��0�E�E;Et�EP�M�E����_^[���   ;���v����]������������������������������U����   SVW��4����3   ������EP�7�����E��}��u2���
�E�M���_^[���   ;��lv����]��������������������������U����   SVW��<����1   ������EP�MQ�S7�������tǅ<���   �
ǅ<���    ��<���_^[���   ;���u����]�����������������������������U����   SVW��4����3   ������E�M���ER��P����B���XZ_^[��]ÍI    ������   ��_Cat �����������������������������������U����   SVW��4����3   ������E�M���ER��P�����XZ_^[��]ÍI    �����   (�_Cat �����������������������������������U����   SVW��4����3   ������E�M���ER��P����B���XZ_^[��]ÍI    ������   ��_Cat �����������������������������������U����   SVW��4����3   ������E�R��P���ʇ��XZ_^[��]ÍI    �����    �_Cat ���������������������������U����   SVW��4����3   ������E�R��P�|��Z���XZ_^[��]ÍI    ������   ��_Cat ���������������������������U����   SVW��@����0   ������E�M��E_^[��]�����������������U���   SVWQ�� ����@   ������Y���3ŉE��M�E�P�M��H���E�P�M Q���̍UR�c�����̍EP�sc���9H���� ������M��j���M��j�������R��P����J���XZ_^[�M�3���V����   ;��r����]� ��   ������   ��_Alval �����������������������������������������������������������������U����   SVWQ��$����7   ������Y���3ŉE��M�E�P�M��G���E�P�MQ�UR�EP�q����R��P����j���XZ_^[�M�3���U�����   ;��q����]� ��   ������   ��_Alval �������������������������������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��4����3   ������M訄����8����M��h����8���_^[���   ;���p����]�����������������������������������U����   SVW��<����1   ������EP�M�R��`�������tǅ<���   �
ǅ<���    ��<���_^[���   ;��=p����]���������������������������U����   SVW��4����3   ������EP�MQ�MX������;�����;���R�EP�MQ�UR�EP��0����_^[���   ;��o����]�����������������������������������������U��j�h0�d�    PQ���   SVW��$����3   �����󫡀�3�P�E�d�    �e�ht  h�]�EP�MQ�Y4����hu  h�]�EP�r�����E�E��E�    ��E��0�E�M��0�M�E;Et�EP�MQ�M��~�����0�	�E��0�E�E�;Et�E�P�M��<����j j �7g���w���E�������E������E�M�d�    Y_^[���   ;��n����]���������������������������������������������������������������������������������U����   SVW��4����3   ������EP�MQ�"_������;�����;���R�EP�w����P�MQ�UR�EP�MQ�Dx����_^[���   ;��m����]��������������������������������������������U��j�h`�d�    PQ���   SVW��$����3   �����󫡀�3�P�E�d�    �e�h�  h�]�EP�MQ�d;����h�  h�]�EP�p�����E�E��E�    ��E��0�E�M��0�M�E;Et�EP�MQ�M��U�����0�	�E��0�E�E�;Et�E�P�M��:����j j �7e���w���E�������E������E�M�d�    Y_^[���   ;��l����]���������������������������������������������������������������������������������U����   SVW������9   ������E$P�M Q��O����P���̍UR�\����x����P���̍EP�|\����x����P�U����P�M Q�g������� ����M��c���M��c���� ���_^[���   ;��k����]���������������������������������������������U����   SVW��@����0   ������EP�MQ� O����P�UR��N����P�EP��N����P��P����P�MQ�Yf����� _^[���   ;���j����]���������������������������������������������U����   SVW��@����0   ������3�_^[��]����������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVWQ��4����3   ������Y�M��EP�A����P�MQ�U�R�W]����_^[���   ;��i����]� ��������������������������U����   SVWQ��$����7   ������Y�M��EPj��M������,�����,��� t$�MQ�~������,���� ���,�����$����
ǅ$���    _^[���   ;��!i����]� ��������������������������������������������U����   SVW��@����0   ������EP�&~����P�MQ�M��K��_^[���   ;��h����]����������������������U����   SVWQ��4����3   ������Y�M��EP�?2����P�MQ�U�R��+����_^[���   ;��?h����]� ��������������������������U����   SVWQ��$����7   ������Y�M��EPj�DL������,�����,��� t*�MQ�1������@��,�����A��,�����$����
ǅ$���    _^[���   ;��g����]� ��������������������������������������U����   SVW��@����0   ������EP�$1����P�MQ�M�/M��_^[���   ;��(g����]����������������������U����   SVWQ��4����3   ������Y�M��EP�S����P�MQ�U�R�LG����_^[���   ;��f����]� ��������������������������U����   SVW��@����0   ������EP�R����P�MQ�M�>��_^[���   ;��Xf����]����������������������U����   SVWQ��4����3   ������Y�M��EP�x.����P�MQ�U�R��q����_^[���   ;���e����]� ��������������������������U����   SVWQ��$����7   ������Y�M��EPj0��I������,�����,��� t)�MQ��-�����   ����,���󥋕,�����$����
ǅ$���    _^[���   ;��Le����]� ���������������������������������������U����   SVW��@����0   ������EP�]-����P�MQ�M��b��_^[���   ;���d����]����������������������U����   SVWQ��4����3   ������Y�M��EP�M�Q�;����_^[���   ;��|d����]� �����������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVW��@����0   ������EP�M�8]��_^[���   ;���c����]�������������������U����   SVWQ��4����3   ������Y�M��EP�M�Q�>����_^[���   ;��c����]� �����������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVW��@����0   ������EP�M�lQ��_^[���   ;���b����]�������������������U����   SVWQ��4����3   ������Y�M��EP�M�Q��B����_^[���   ;��b����]� �����������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVW��@����0   ������EP�M�N��_^[���   ;��b����]�������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������E_^[��]�������������������������U���   SVW�������H   �����󫡀�3ŉE�j �M��82������E����\.���E܋E�P�M�U���EЃ}� t�|�}� t�E�E��n�EP�M�Q�I�������u#h|]�������L7��hH=������P�X���6�E�EЋE����E�EċEċ��MċB��;���_���E�P�c�����EЉ������M���\��������R��P�� 	�Zs��XZ_^[�M�3���C����   ;��_����]�   � 	����   � 	����   � 	_Psave _Lock �����������������������������������������������������������������������������������U���   SVW�������H   �����󫡀�3ŉE�j �M��0������E蹈��,���E܋E�P�M�T���EЃ}� t�|�}� t�E�E��n�EP�M�Q�jX�������u#h|]�������5��hH=������P��V���6�E�EЋE����E�EċEċ��MċB��;��A^���E�P�qa�����EЉ������M��1[��������R��P�0	�q��XZ_^[�M�3��:B����   ;���]����]�   8	����   W	����   P	_Psave _Lock �����������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���U���M���E�_^[���   ;��/]����]�����������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@   �M��R���E�_^[���   ;��\����]����������������������������U����   SVWQ��4����3   ������Y�M��M���_���E�_^[���   ;��a\����]�������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��J���E�_^[���   ;���[����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��_���E�_^[���   ;��[����]�������������������������������U����   SVWQ��4����3   ������Y�M��M��3���M��F���E�_^[���   ;��9[����]� ��������������������U����   SVWQ��4����3   ������Y�M��M��W���EP�M��Y���E��M�H�E�_^[���   ;���Z����]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M��a%���E�_^[���   ;��iZ����]� ��������������������U����   SVWQ��4����3   ������Y�M��M��4T���E��@    �E��@    �E�_^[���   ;���Y����]���������������������������U����   SVWQ��4����3   ������Y�M��M��jg���M��Y*���E�_^[���   ;��Y����]� ��������������������U����   SVWQ��4����3   ������Y�M��EP�M��(���E��M�Q�P�E�_^[���   ;��1Y����]� ����������������������������U����   SVWQ��4����3   ������Y�M��M��$���E��M�H�EP�M��W���E�_^[���   ;��X����]� �����������������������U����   SVWQ��4����3   ������Y�M��M��R���E��@    �E��@    �E��@    �E�_^[���   ;��CX����]���������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��;���E�_^[���   ;���W����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��9b���E�_^[���   ;��W����]�������������������������������U����   SVWQ��4����3   ������Y�M��M���1���E�_^[���   ;��!W����]�������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��%>���E�_^[���   ;��V����]� ������������������������U����   SVWQ��4����3   ������Y�M��M���,���E�_^[���   ;��aV����]�������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@ �E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��E��     3��M�f�A�E�_^[��]������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��M���V���E�� LUj �EP�M���#���E�_^[���   ;��
T����]� �������������������������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �} t�E�� �U�M���p�����,���j j �E���P�M��;���E���Q�E���U�E���Q��p�E���A�M��T�j �M�����<���EP�M��Q�UR�M����(����uj j�E���U�Q���e���E�_^[���   ;���R����]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��"���E�� �T�E�_^[���   ;��xR����]����������������������U����   SVWQ��(����6   ������Y�M�ǅ,���    �} t�E�� �T�M��������,����E���Q�E���T�E���Q���E���A�M��T��E��@    �@    �EP�MQ�U���M�H�2?���E�_^[���   ;��Q����]� ���������������������������������������������������U����   SVWQ��$����7   ������Y�M��E��  Ujh�[��J��Pj�*e������,�����,��� t��,����\����$����
ǅ$���    �E���$����H4�M���7���E�_^[���   ;���P����]���������������������������������������U����   SVWQ��(����6   ������Y�M���/���P�M��T��P�M�����j j �M��&���EP�~O����P�M������E�_^[���   ;��@P����]� �������������������������������������������U����   SVWQ������9   ������Y�M���/���P��#���Q�M�@T�����S��P�M��9��j j �M��g%���@QPj �MQ�M��O���E�_^[���   ;��O����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M���/�����Y��P�M����j j �M���$���EP�MQ�M��JG���E�_^[���   ;���N����]� �����������������������������������U����   SVWQ��(����6   ������Y�M���/����FY��P�M����j j �M��9$���EP�M������E�_^[���   ;��mN����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M���/����X��P�M��{��j j �M��#���E�_^[���   ;���M����]�����������������������U����   SVWQ��4����3   ������Y�M��EP�M��b'���E�� �Z�EP�M������E�_^[���   ;��xM����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��;���E�� �R�EP�M���>���E�_^[���   ;���L����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E��     �@    �E��M�H�U�P�E��M�H�E�_^[��]� �������������������������U����   SVWQ��4����3   ������Y�M��E��M��U�P�E��@    �@    �E��@    �E�_^[��]� ������������������������U��j�h��d�    PQ���   SVWQ�������?   ������Y���3�P�E�d�    �e��M荅���P������Q�M�Y!������E��P�M��%���M�2X��P�M���F������t]�E�    �E�HQ��T�M�#����T�M�M/���M������U�B��M���"��j j �C���
	��E�������E������E�M�d�    Y_^[��  ;���J����]� ���������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M���/����� ��P�M��u$���E�_^[���   ;��UJ����]�����������������������������������U����   SVWQ��4����3   ������Y�M��E��M��E��M�H�E��M�H�U��E�B�E�_^[��]� ������������������������������U����   SVWQ��4����3   ������Y�M��M���2���E�� ,P�E�_^[���   ;��xI����]����������������������U����   SVWQ��4����3   ������Y�M��E��E� �E��E�@�E��E�@�E�_^[��]� ���������������������������U����   SVWQ��4����3   ������Y�M��E��x^� �E��x^�@�E��x^�@�E�_^[��]�������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E��@    �E��@    �E��@    �E�_^[��]�������������������������������U����   SVWQ��4����3   ������Y�M��M��A3���E�� �U�E�_^[���   ;��G����]����������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��>G����EPj��MQ�U�R����H�Q�҃�;��G���E�_^[���   ;��G����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��F���E�_^[���   ;��{F����]�������������������������U����   SVWQ��4����3   ������Y�M��E��     �E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E�� lQ�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��M��L=���E�� XS�E�_^[���   ;��(E����]����������������������U����   SVWQ��4����3   ������Y�M��M������E�� �S�E�_^[���   ;���D����]����������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �EP�M���%���E�_^[���   ;��ZD����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVWQ�� ����8   ������Y�M�j �M��m���M����A���M����A���M����O���M����O���M���$��@���M���,��@���} u!hTQ��$����#��hT<��$���P��;���EP�M�Q�������E�_^[���   ;��&C����]� �������������������������������������������������U����   SVWQ��,����5   ������Y�M��E��M��E����0�����0������0���H�����tC�E����0�����0������0���H�e����,�����,������,����B��;��\B���E�_^[���   ;��IB����]� ����������������������������������������������������U����   SVWQ��,����5   ������Y�M��E��M��E����0�����0������0���H�����tC�E����0�����0������0���H�����,�����,������,����B��;��|A���E�_^[���   ;��iA����]� ����������������������������������������������������U����   SVWQ������?   ������Y�M����̋EP����MQ�UR�����P������(P�M���T��������A���E�� 4S�E��M�H�U�P�E�_^[���   ;��@����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��j&���E�� 4S�E�H�P�E��H�P�E�_^[���   ;��"@����]� �����������������������������U����   SVWQ��4����3   ������Y�M��M�����E�� �S�E�_^[���   ;��?����]����������������������U����   SVWQ��4����3   ������Y�M��EP�M��� ���E�� �Q�E�_^[���   ;��T?����]� �������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��o ���E�� �R�E�_^[���   ;���>����]� �������������������������������U����   SVWQ��4����3   ������Y�M��E�� S�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E��M��E��M�H�E�_^[��]� ����������������U����   SVWQ��4����3   ������Y�M��E��M��E��M�H�E�_^[��]� ����������������U����   SVWQ��4����3   ������Y�M��M��A ���E�� �Q�EP�M���Q������E�_^[���   ;��u=����]� ��������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��x&���E�� T�E�_^[���   ;��=����]� �������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�QR�P�M��[7���E�� T�E�_^[���   ;��<����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��E�_^[��]� �������������������������U����   SVWQ��4����3   ������Y�M��E��  T�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E��M���E���U����
�P��;��x;���E�_^[���   ;��e;����]� ��������������������������������U����   SVWQ��4����3   ������Y�M�j�e,�����M���E�_^[���   ;���:����]������������������������U����   SVWQ��4����3   ������Y�M��E��E� �E��E�@�E��E�@�E�_^[��]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�M���B���E�� HQ�E�_^[���   ;��$:����]� �������������������������������U����   SVWQ��(����6   ������Y�M��M�/����,�����,���P�M��Z���E�� HQ�E�_^[���   ;��9����]� ������������������������������U����   SVWQ��4����3   ������Y�M��EP�M������E�� HQ�E�_^[���   ;��49����]� �������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��Z���EP�M��	��H���U��B�E�_^[���   ;��8����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�����E��UQ���Q�������tF�E��UQ���"(����t0�E��UQ���(��;Et�E��UQ����'�����3���E��UQ��������M��A�E�_^[���   ;���7����]� �������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M�����E��P�M�������E�_^[���   ;��K7����]� ����������������������U����   SVWQ��4����3   ������Y�M��EP�M��!���M��������M�[
���E�_^[���   ;���6����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��b���E�� HS�E�_^[���   ;��d6����]� �������������������������������U����   SVWQ������<   ������Y�M��EP������=�������Q�UR�EP�M����������Y	���E�� HS�E�_^[���   ;���5����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��U�P�M�H�E����M��U�P�M�H�E����M,��U0�P�M4�H�E���$�M ��U$�P�M(�H�E�_^[��]�0 ����������������������������������������U����   SVWQ��4����3   ������Y�M��E�P�������E��     _^[���   ;��4����]���������������������U����   SVWQ��4����3   ������Y�M��M��)��_^[���   ;��T4����]������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;��4����]������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;��3����]������������������U����   SVWQ��4����3   ������Y�M��M��L)���M��D��_^[���   ;��\3����]��������������������������U����   SVWQ��4����3   ������Y�M��M��;��_^[���   ;��3����]������������������U����   SVWQ��4����3   ������Y�M��M��!���_^[���   ;��2����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��d2����]������������������U����   SVWQ��4����3   ������Y�M��M������M������_^[���   ;��2����]��������������������������U����   SVWQ��4����3   ������Y�M��M��J���_^[���   ;��1����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��d1����]������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;��1����]������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;���0����]������������������U����   SVWQ��4����3   ������Y�M��E�� LU�E��xP t�M�����E��HL��t�M��j ���M������_^[���   ;��G0����]�������������������������������������U����   SVWQ��4����3   ������Y�M��E��H��Q�E��D��U�E��H��Q��p�E��H��A�M��T��M���`�>���M���X����_^[���   ;��/����]������������������������������������U����   SVWQ��4����3   ������Y�M��E�� �T�M����_^[���   ;��;/����]�������������������������U����   SVWQ��4����3   ������Y�M��E��H�Q�E��D��T�E��H�Q���E��H�A�M��T�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��E��  U�E��H4Q�>�����_^[���   ;��d.����]����������������������������������U����   SVWQ��4����3   ������Y�M�j j�M�����M��#��_^[���   ;���-����]����������������������U����   SVWQ��4����3   ������Y�M��E�� �Z�M��Q��_^[���   ;��-����]�������������������������U����   SVWQ��4����3   ������Y�M��E�� �R�M��2#���M�����_^[���   ;��3-����]���������������������������������U����   SVWQ��4����3   ������Y�M��M�����M������_^[���   ;���,����]��������������������������U����   SVWQ��4����3   ������Y�M��M��7��_^[���   ;��t,����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��$,����]������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;���+��_^[���   ;��+����]����������������������������U����   SVWQ��4����3   ������Y�M��M��j��_^[���   ;��d+����]������������������U����   SVWQ��4����3   ������Y�M��E�� lQ_^[��]��������������U����   SVWQ��4����3   ������Y�M��M��y��_^[���   ;���*����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��*����]������������������U����   SVWQ��$����7   ������Y���3ŉE��M�j�M�������M��a���M��5'��R��P�(6	��=��XZ_^[�M�3��D�����   ;���)����]Ë�   06	����   <6	_Lock ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E�P�-�����M���,�i+���M���$�^+���M����j���M����_���M����=+���M����2+���M��C&��_^[���   ;��&)����]������������������������������������U����   SVWQ��,����5   ������Y�M��E����0�����0������0���H������tC�E����0�����0������0���H�}�����,�����,������,����B��;��t(��_^[���   ;��d(����]��������������������������������������������������U����   SVWQ��,����5   ������Y�M��E����0�����0������0���H�������tC�E����0�����0������0���H������,�����,������,����B��;��'��_^[���   ;��'����]��������������������������������������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��$'����]������������������U����   SVWQ��4����3   ������Y�M��M������_^[���   ;���&����]������������������U����   SVWQ��4����3   ������Y�M��E�� �Q�M�����_^[���   ;��{&����]�������������������������U����   SVWQ��4����3   ������Y�M��E�� �R�M��&���_^[���   ;��&����]�������������������������U����   SVWQ��4����3   ������Y�M��E�� S_^[��]��������������U����   SVWQ��4����3   ������Y�M��E�� �Q�M��]��_^[���   ;��{%����]�������������������������U����   SVWQ��4����3   ������Y�M��M��{��_^[���   ;��$%����]������������������U����   SVWQ��4����3   ������Y�M��E��  T�E�P������_^[���   ;���$����]���������������������U����   SVWQ��4����3   ������Y�M��E��8 t#�E���U����
�P��;��j$��P�������_^[���   ;��Q$����]�������������������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;���#����]������������������U����   SVWQ��4����3   ������Y�M��M���7��_^[���   ;��#����]������������������U����   SVWQ��4����3   ������Y�M��������u
�E���/���M�����_^[���   ;��>#����]����������������������������U����   SVWQ��4����3   ������Y�M��M����:����M��W���_^[���   ;���"����]�����������������������U����   SVWQ��4����3   ������Y�M��M��O���_^[���   ;��"����]������������������U����   SVW��@����0   ������E_^[��]�������������������������U����   SVW��@����0   ������EP�MQ�UR�EP��5����_^[���   ;���!����]�����������������������U����   SVW��@����0   ������EP�"�����_^[���   ;��!����]�������������������U����   SVWQ��$����7   ������Y���3ŉE��M�E�M�;u�4�E�8 t�E��R�M������j�M�������M��I����M�����E�R��P�D?	�4��XZ_^[�M�3��)�����   ;��� ����]� �   L?	����   X?	_Lock ��������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��u��_^[���   ;��T ����]������������������U����   SVWQ��0����4   ������Y�M��E�;Euǅ0���   �
ǅ0���    ��0���_^[��]� ��������������������������������U����   SVWQ��0����4   ������Y�M��M�9��P�M��0������������t"�M�������M���;�uǅ0���   �
ǅ0���    ��0���_^[���   ;��K����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|.h�Zh�   h�ZhL[������h�Zh�   �J0����kE�M�A_^[���   ;������]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M��M���*��;Ewhh�  h0Xh�X�e����� Y��t3�u&hPYh�Yj h�  h0Xj�k�������u�j h�  h0Xh�Yh�Z�"����kE0�M�A_^[���   ;������]� ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M��Q�pq��_^[��]������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��$����7   ������Y���3ŉE��M�E�8 u2j �M��k����E�8 u�|����|��M�|���M�����E� R��P��C	�0��XZ_^[�M�3�� �����   ;��X����]Ð   �C	����   �C	_Lock ����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��M�������tD�E��x t;�M�����������M�9Ar$�M��r�����������M��a���p�E�;pw_jOh�Vh \������� Y��t3�u#hPYh�Yj jPh�Vj���������u�j jPh�VhX\h�Z������E��@_^[���   ;��W����]���������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;�������]������������������U����   SVWQ��4����3   ������Y�M�j�j��EP�M��W&��P�M�����E�_^[���   ;��p����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M���p�u)���M���p���_^[���   ;������]��������������������U����   SVWQ��4����3   ������Y�M��M���������M����\��_^[���   ;������]��������������������+I��w����+I��9����������������U����   SVWQ��4����3   ������Y�M��M��&���E��t�E�P�,�����E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M���p����E��t�E���pP�+�����E���p_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�+�����E�_^[���   ;��-����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��������E��t�E���P�*�����E���_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�!*�����E�_^[���   ;��=����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��P����E��t�E�P�������E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M��3*���E��t�E�P�5������E�_^[���   ;��]����]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P��(�����E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�a(�����E�_^[���   ;��}����]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P��'�����E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�'�����E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�'�����E�_^[���   ;��-����]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�&�����E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M��_'���E��t�E�P�1&�����E�_^[���   ;��M����]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�������E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�E������E�_^[���   ;��m����]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P��$�����E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�e������E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�$�����E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�#�����E�_^[���   ;������]� ������������������������U����   SVWQ��4����3   ������Y�M��M��W����E��t�E�P�!#�����E�_^[���   ;��=����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��E����E��t�E�P�"�����E�_^[���   ;�������]� ������������������������U����   SVWQ��4����3   ������Y�M��M�������E��t�E�P�A"�����E�_^[���   ;��]����]� ������������������������U���h  SVWQ�������  ������Y���3ŉE��M�j�M�������M������j h�U�������������������P������Pj j�M�� ������������������������j hV�����������������P�M���������������������������� �4  j�M��#����M������h1D4ChCD4Cjjj�E�P�M���������[�����u%ǅ����    �M������M�������������  j�M��u��j h�Q�M��1����M��������Z����E�ǅ ���   �� ���s������ ����D� �   k� �T��U�ǅ|���    ���|�������|�����|���;E�tE�E�P�M��$����������j �E�P���������P�M����������w�����|���~��j hV��$����n���j j ��$���P�M��6�����t	ƅ�����ƅ���� ��������s�����$��������M�������������s������`  j ��<���P�M���������#��P�������^��������Q��<���R������������������<��������M��e��j��$���������$���P�M�����j������������X���P������{�������������� ���k� ����������� ���Pk� ���Q����������������������������������"�������������������������������p����u���j��P����i�����P����Q���ǅD���    ���D�������D�����D���;������~  k�D�����8���k�D�������,���k�D������� �����D���;� �����  ��D���P����������Z@���$��D���Q������g����Z@���$��D���R������H����Z@���$��T����%�����������P�������H�������P�������H�������P��������D���P�����������Z@ ���$��D���Q�����������Z@���$��D���R����������Z@���$��t���������������P�������H�������P�������H�������P��������D���P������L����Z@,���$��D���Q������-����Z@(���$��D���R����������Z@$���$��������������p����P��t����H��x����P��|����H�������P���������ċ�������������P�������H�������P�������H�������P��P�����������ċ�������������P�������H�������P�������H�������P��P����������ċ�p������t����P��x����H��|����P�������H�������P��P����H�����D���;� ���}E�� ���P��,���Q��8���R������������D�������������P�Q�P�Q�@�A��D���P��P�������k�D�����������P�Q�P�Q�P�Q�P�Q�@�A�a���j j�������$���j j j ������P�M�����j����������������&����������4����E�����������������������������jh  ���������jh  �������������^�$h  ��������������Ph�   �e�����ǅ����    ��X����*����<����L���E�    �E�P�������E�������������Q������������ uǅ����    ��E�#�  �U�������j ��P����2�����P������������������������������P����>��������������$���������<����	����.j hV����������j0������P�������������n����M��f����M�����j ������ǅ����   �M�����������R��P�,[	����XZ_^[�M�3��@�����h  ;�������]�    4[	����   "\	����   \	����   \	����   \	����   \	<���,   \	$���   \	���   \	����   �[	����   �[	p���   �[	P���   �[	���   �[	����   �[	mdat bc tri_positions posc posb posa triangles name info pc c text bf file �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M��B@��;����_^[���   ;������]� ����������������������������������U����   SVWQ������9   ������Y�M��E��8 tD�E�    �E��H�M��E�    ��E���E�M����M��E��M�;H}��E�P��������E��     �E��@    �E��@    �E��@    �E��@    _^[���   ;��/ ����]�������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�����P��M��B<��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M��h���_^[���   ;��=�����]���������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M�����_^[���   ;��������]���������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���   �҃�;��t���_^[���   ;��d�����]� �������������������������������U����   SVWQ��4����3   ������Y�M��}  }3��Njjj�E P�M��������u3��4kE �M��QЋE��M�J�E�B�M�J�E�B�M�J�   _^[���   ;�������]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M��BL��;��2���_^[���   ;��"�����]� �����������������������������U���P  SVWQ�������T   ������Y�M��} }3��  �} 
�   �  �E��H;M~�U��B�������	�M������������U�U�E��x uh�ZhA  �����3��4  �E��H��9M��  �E��H+M�U��J�E��x �s  �E��@�؃��M���y���U��B��E܉U��E��@�E�U�j jRP�|���ẺUЋE̙�������������E�;�����ud�M�;�����uY�E��@�E�U��������������M�;�����|5�U�;�����r(�E��������������E�;�����K|�M�;�����s>�   ��t.h�]hP  h�ZhL[�n�����h�ZhP  ������3��	  �E܋M�A�U��B�E܋M�A�U��B�E��8 u6��h�ZhW  �E�kHQ����B���  �у�;�������U���:��h�ZhX  �E�kHQ�U��P����Q��  �Ѓ�;������M���E��8 u3��d  �E�kH�U�
�E��H�} ~�E��H+Mk�R�E��ȋ�+M�u��E���j jVQ�����U�BP�EEk��U�JQ�B�����kEP�E�+E�U�j jRP����M�AP�U��BP�������7�E�kHQ�E�+E�U�j jRP�`���U�BPkE�M�AP��������9�} ~!kEP�M��QR�E�kH�U�
Q�������E�kH�U�
�E��H��  �E��H�U�D
��M���y���U��B��E��U��E��@��������������M�;������a  �U�;������P  j j�E�P�M�Q����E��U��E���������������E�;�����uE�M�;�����u:�E�;E�|2�M�;M�r(�E��������������E�;�����K|�M�;�����s>�   ��t.h�]hx  h�ZhL[������h�Zhx  �
����3��I  �E��8 u3��h�Zh|  kE�P����Q���  �Ѓ�;��P����M���6��h�Zh}  kE�P�M��R����H��  �҃�;������M���E��8 u3���  �E�kH�U�
�E��H�E��M��A�E��M;H}0�E��H+Mk�RkE�M�AP�UUk��M�AP�������E�    �E�    �} t_�E��H;M}1�E�kH�U�JQ�E��M+Hk�R�E�kH�U�JQ�������kE�M�APkURkE�M�AP�������} ��   �E��H;M}q�E��H�M��U�kB�M�A�E���E����E��M����M��E�;E}<�E�Pj�9����������������� t�������k����������
ǅ����    ��E�    kE�M�A�E���E����E��M����M��E�;E}<�E�Pj������������������� t������������������
ǅ����    몋E��M�H�   _^[��P  ;��+�����]� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ������   �M��P��;��'���_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��HQ���ԋE��M�J�E�B�M�J�E�B�M�J�M��5��_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M��E��M;Hu�   �@�E��M;H}�E��H+MQ�UR�M��,����jj�E��M+HQ�U��BP�M��ɾ��_^[���   ;��������]� �������������������������������������U���  SVW�������F   ������hHV� ���Ph��j������������������ t�����������������
ǅ����    j h�V��,����d���������Qj h�V������K���P��,���R�� ��������������Pj h'  ������Ph�� �������������� �������������������,��������������_^[��  ;�������]����������������������������������������������������������������������U���  SVWQ�������E   ������Y�M��} 
�   ��  �} |�E��M;H}�E��8 u3��  �E��x uh�Zh�  �~����3��  �} �E��M;H|�M������   �q  �E��HQ�UUR��������E�E�+E�E��E�    �E�    �E�    kE�M�A�E���Eԃ��EԋMȃ��MȋE�;E�}��E��H��9M�  �E��HM��U��J�} ~kEP�M��QRkE��M�AP�(������E�kH�U�
�E��H�E��M��P;Q��   �E��M��@��y�U��B�E��E��H+M��U��J�E��H+M��U��J�E��H+M�k�R�E��HQ�U���k��M�AP褽������h�Zh�  �E�kHQ�U��P����Q��  �Ѓ�;��g����M���E��8 u3���   �E�kH�U�
�E��H��   �E��H�U��B�D�+E��M���y���U��B�E��E��H��9M}5�EE��M��Q+�k�P�MM�k��E�PRkM�U�JQ�ڼ�����E��M�;H}]��h�Zh�  kE�P�M��R����H��  �҃�;������M���E��8 u3��/�E�kH�U�
�E��H�E��M��H�E��H+M��U��J�   _^[��  ;��F�����]� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��P0��;��*���_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�EP����Q�M��B,��;�����_^[���   ;�������]� ����������������������������U����   SVW��@����0   ������E;E}�E��E_^[��]����������������������������U����   SVWQ������=   ������Y���3ŉE��M�} uj�M�蝽���M������M�������I�E��M܋E�;M�t7j�M��o����M�������E�M܋Q�P�E܋M�H�E�M܉�M�����R��P��t	�#���XZ_^[�M�3��������   ;��\�����]� �I    �t	����   �t	����   �t	_Lock _Lock ������������������������������������������������������������������������U����   SVWQ������;   ������Y���3ŉE��M�M��u���j�M��v����M����������P�E�Q�M��x����E��U�R��P��u	����XZ_^[�M�3��������   ;��L�����]Ð   �u	����   �u	_Alproxy �����������������������������������������������������������U����   SVWQ������;   ������Y���3ŉE��M�M�����j�M��y����M����������P�E�Q�M������E��U�R��P��v	�#���XZ_^[�M�3��������   ;��\�����]Ð   �v	����   �v	_Alproxy �����������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�xs"�E�H��Q�U��R�E���P�s������.�E��P�M���Q��/���R�M���������~����E�@    �E��M�Q�P�E��M�Q�Pj j �M����_^[���   ;��O�����]� ����������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��@    �E��@    �E��@    �} u2��W�S�M�����;Es
�M������<�EP��/���Q�M��^������}����U��B�E��M��Q�PkE0�M�A�U��B�_^[���   ;��]�����]� ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M��}u�EP�M�����EP�+�������EP�MQ�M�����EP������_^[���   ;�������]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     _^[��]��������������U��j�h��d�    PQ��  SVWQ�������C   ������Y���3ŉE�P�E�d�    �e��M�E���E؋M��d���;E�s�E�E��R�E�H��E�3Ҿ   ��;�w�8�M��5����M�Q��+M�9Aw�E�H��U�J�M���M������E��E�    �E؃�P������Q�M��������輮���E��`�e��E�E��E��E؃�P������Q�M�������荮���E��j j�M��Ϻ��j j �����{	��E�   ��E�   �+{	��E�������E������} v�EP�M�����P�M�Q�m�����j j�M��o����E�P�M��Q�����R�M�������蒭���E�M؉H�EP�M������R��P��{	�(���XZ�M�d�    Y_^[�M�3�������  ;��V�����]� �   �{	����   �{	_Ptr ���������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��������Iu�E���3�_^[��]������������������������������U����   SVWQ��$����7   ������Y���3ŉE��M�E�P�M��ܸ���E�P�MQ�UR�������R��P�P}	����XZ_^[�M�3��������   ;��������]� ��   X}	����   d}	_Alval �����������������������������������������������������U����  SVWQ��(����v   ������Y���3ŉE��M�ǅ����    �E�x@ t�E��HE��u��E  �@  �E�   �������P�E��M�B��;�������0���������<�����0���Q��<���R�����������t2���  j j�M��Ĺ���E�P��T���Q�M��������������M������V��h���R�M�����������P�E��HP�M�I@������H�����h���������T���������H�����(�����(��� t��(���t��(����
  �  �E��@E ��|���P�M������������M�+ȉM���|����D����}� vD�E�HPQ�U�Rj������P�M�������������������P�������9E�tǅ(���   �
ǅ(���    ��(�����������������t��������������������������tƅ���� �M��ϳ���������q�E��HE��uƅ�����M�譳���������O�}� uj j�M�萻���.ƅ�����M�肳���������$ƅ���� �M��k�����������,����M��V���R��P�h�	����XZ_^[�M�3��������  ;�������]Ë�   p�	����   ��	����   ��	_Str _Dest ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�ƅ/��� �E��M�H��/���R�M��F���EP�������_^[���   ;��q�����]� ����������������������������U����   SVWQ��$����7   ������Y���3ŉE��M�M������M������E�Q�M��k���j�E�Q�M������E��     R��P�d�	����XZ_^[�M�3��������   ;��������]Ð   l�	����   x�	_Alproxy �����������������������������������������������U����   SVWQ��$����7   ������Y���3ŉE��M�M�蝬���M��(����E�Q�M�����j�E�Q�M��"����E��     R��P�D�	����XZ_^[�M�3��'������   ;��������]Ð   L�	����   X�	_Alproxy �����������������������������������������������U����   SVW��@����0   �������EP�MQ����B��0  �у�;��L���_^[���   ;��<�����]��������������������������U����   SVWQ��4����3   ������Y�M��M�m����E_^[���   ;��������]� ����������������������������U����   SVWQ��4����3   ������Y�M��M�����E_^[���   ;�������]� ����������������������������U���  SVW�������F   ������ǅ8���    �} ��   �E�8 ��   h�  h�Q�����Pj�I����������������� t1j �M�����P�������]�����8���P������������������
ǅ����    �E���������8�����t��8���������������   _^[��  ;�������]��������������������������������������������������������������U���  SVW�������F   ������ǅ8���    �} ��   �E�8 ��   h�	  h�Q����Pj�)����������������� t1j �M����P�������=�����8���P������藵���������
ǅ����    �E���������8�����t��8�����������f����   _^[��  ;��`�����]��������������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��8 uǅ0���    ��M�����0�����0���_^[��]��������������������������������U����   SVWQ������?   ������Y�M��� ���P�������������P������H������P������E������������P������H������P�E_^[���   ;��!�����]� ��������������������������������������������U����   SVWQ������:   ������Y�M��E���U;Qs�E���Q�E��������
ǅ���    ������U�}� u�E���Q��u�E��9�7������E��E��M;Hs�U��B�M��������
ǅ���    �����_^[���   ;��5�����]� ������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��8 uǅ0���    ��M������0�����0���_^[��]�������������������������������U����   SVWQ��4����3   ������Y�M��E���_^[��]�����������������U����   SVWQ��0����4   ������Y�M��E��H�9 t�U��B,���0����
ǅ0���    ��0����_^[��]���������������������������U����   SVWQ��0����4   ������Y�M��E��H,����E��H,��E��H�����0����E��H��0������0���_^[��]�������������������������������U����   SVWQ��0����4   ������Y�M��E��H,����E��H,��E��H���0����E��H����E��H���0���_^[��]�����������������������������U����   SVWQ��0����4   ������Y�M��E��H,����E��H,��E��H�����0����E��H��0������0���_^[��]�������������������������������U����   SVWQ��0����4   ������Y�M��M�����;Es�M�肿���E��H;Ms�E��HQ�UR�M������S�E��t;�}s5�E��M;Hs�U��0�����E��H��0�����0���Rj�M��s�����} u
j �M�� ����} vǅ0���   �
ǅ0���    ��0���_^[���   ;�������]� �������������������������������������������������������������U����   SVWQ��$����7   ������Y�M��M�������E�M��[����M���+�;E�sǅ$���    ��U���U쉕$�����$����E�E�;Es�E�E�E�_^[���   ;�������]� ������������������������������������U����   SVWQ��4����3   ������Y�M��E����   ��_^[��]������������������������U���   SVWQ�� ����@   ������Y�M��}uǅ ���   �
ǅ ���    �E��� ����HL�E��@E �M��۸���} tJ�   ��tA�E���E�E�E��E���EԋE���EȋE�P�M�Q�U�R�E�P�M�Q�U�R�M������E��M�HP�E�����HH�E��@@    _^[��   ;��f�����]� �����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M�H�E��M�H�E��M�H�E��M�H �E��M�H,�E��M�H0_^[��]� ������������������������������U����   SVWQ��4����3   ������Y�M��E����M��A�E����M��A�E����M��A�E����M��A �E���$�M��A,�E���(�M��A0j j �M��Ե��j j j �M������_^[���   ;��
�����]����������������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ������9   ������Y�M��� ���P�M诒���M������P�Q�P�Q�@�A_^[���   ;��A�����]� ����������������������������U����   SVWQ��$����7   ������Y�M��E��@0    �E��@    �E��@    �E��@  �E��@   �@    �E��@     �@$    �E��@(    �E��@,    j �M��l���h  h�T�E���Pj�x�������,�����,��� t��,����������$����
ǅ$���    �E���$����H0_^[���   ;��2�����]����������������������������������������������������������������U����   SVW��@����0   ������E�M�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��M�ӗ������t�E��@@    ��E��M�H@�M��V���_^[���   ;��P�����]� ���������������������������U����   SVWQ��4����3   ������Y�M��} t �M�跴��9Er�M�誴���M�A;Ew2����_^[���   ;��������]� �������������������������U����   SVWQ��0����4   ������Y�M��E��M;Hs�U��B;Ewǅ0���   �
ǅ0���    ��0���_^[��]� ����������������������������������U��j�h �d�    PQ��   SVWQ�������@   ������Y���3ŉE�P�E�d�    �e��M�E��U�Q���׌�������t  �E��U�Q��褻����t�E��U�Q��莻�����D����E���  �E��U�Q����������  ������P�M��M�J�_���P�������E؍������8����E�    �E��U�Q��������������E���E��U�Q����������t����E������� ����E�P�� ���Q�ݸ�����Ѕ�tj j�E��U�Q��������'�#�E�P���������QjH�M�������Ѕ�u���jj�E��U�Q���������	��E�������E������E��U�Q���c�������t��j j�E��U�Q���F���2�R��P� �	�����XZ�M�d�    Y_^[�M�3��N�����  ;�������]� ��   (�	����   4�	_Meta ������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��xP t�E��HPQ�������_^[���   ;�������]����������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVW������9   ������M���������uh@S�M�p����� ���P�M����P�M�߮���� ���谛���EP�M�;����M蜛���E_^[���   ;�������]�����������������������������������������U����   SVWQ��0����4   ������Y�M��E��xr�M��QR藵������0�����E�����0�����0���_^[���   ;�������]����������������������������������������U����   SVWQ��0����4   ������Y�M��E��xr�M��QR��������0�����E�����0�����0���_^[���   ;��������]����������������������������������������U����   SVWQ������:   ������Y���3ŉE��M�E�8 tMj�M��K����E����M���E܋�U܋A��E܃8 t�E܋�    �ދE��A    �M��Z���R��P��	�����XZ_^[�M�3��i������   ;��"�����]ÍI    �	����   �	_Lock ������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��8 t]�E�����M�E�8 t�E�;M�t�E����M���E�8 uh�   hXPhQ舮�����E�M��Q��E��     _^[���   ;��'�����]�����������������������������������������������������U����   SVWQ������:   ������Y���3ŉE��M�j�M��s����M�贶���E܃}� tN�E܃8 tF�E܋�Q;Ur�E܋�U;Qs�E܋�)����E���E܋������E܋�����M܋�벍M��^���R��P� �	�����XZ_^[�M�3��m������   ;��&�����]� �   �	����   �	_Lock ����������������������������������������������������������������������U��j�h@�d�    PQ���   SVWQ��$����3   ������Y���3�P�E�d�    �e��M��E�    �E��U�Q���c�������tK�E��U�Q��������t4�E��U�Q��������論�����uj j�E��U�Q��������"�	��E�������E������M�d�    Y_^[���   ;��������]�������������������������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��H �9 t�U��B0���0����
ǅ0���    ��0����_^[��]���������������������������U����   SVWQ��0����4   ������Y�M��E��H0����E��H0��E��H ���0����E��H ����E��H ���0���_^[��]�����������������������������U��j�hp�d�    PQ��  SVWQ�������B   ������Y���3�P�E�d�    �e��M�EP������Q�M��������+����E��E�    �E�P�M�QR�E�HQ�M�������-�EP�M�Q������R�M��Ȗ���������j j �r����<�	��E�������E������M������EЋE�x tH�E�HQ�U�BP�M��v����E�M�@+A��0   ��P�U�BP�����Q�M��M������u����M��n���kE0E܋M�AkE�0E܋M�A�E�M܉H�M�d�    Y_^[��  ;��:�����]� �����������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��Q���;Es>�M��������M��D���+�;us�M������M��-���EP�M��l���P�M�����_^[���   ;��Q�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��q����M���D;�u�E��H<Q�U��B8P�M��Q8R�M�誯��_^[���   ;�轾����]���������������������������U����   SVWQ��4����3   ������Y�M��M������M���D;�t�M��ߠ���M��A8�M��c����M��A<�E���EP�M���DQ�U���DR�M�����_^[���   ;��!�����]�����������������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 tj�E��Q�ő�����E��     _^[���   ;�蛽����]�������������������������U����   SVWQ��4����3   ������Y�M��E��8 tj�E��Q�U������E��     _^[���   ;��+�����]�������������������������U����   SVWQ������<   ������Y�M��E��u�y�E��xrp�E��H�M�E���P�����Q�M��$����������} v �EP�M�Q耪����P�U���R�,������E��H��Q�U�R��#���P�M���������6����E��@   �EP�M�迌��_^[���   ;��C�����]� ��������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x ~�E��HQ�X������$�E��x }�E��H��,�����,���R譠�����E��HQ�#�����_^[���   ;�������]���������������������������������������������U����   SVWQ��(����6   ������Y�M��E��x tn�M������E��HQ�U��BP�M��Ɉ���E��M��@+A��0   ��P�U��BP��/���Q�M�蠐������z���E��@    �E��@    �E��@    _^[���   ;�襺����]���������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��xP t�E��HPQ蚼����_^[���   ;�������]����������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��E��M��@+A��0   ��_^[��]�������������������U����   SVWQ��4����3   ������Y�M�h\[�G���_^[���   ;�������]��������������������������������U����   SVWQ��4����3   ������Y�M�h�[�����_^[���   ;�蒸����]��������������������������������U����   SVWQ��4����3   ������Y�M�hp[�B���_^[���   ;��2�����]��������������������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q�_�����_^[���   ;��ʷ����]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q�������_^[���   ;��j�����]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q蟣����_^[���   ;��
�����]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q�?�����_^[���   ;�誶����]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q�ߢ����_^[���   ;��J�����]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q������_^[���   ;�������]� ���������������������U����   SVWQ��4����3   ������Y�M��EPj �M�Q������_^[���   ;�芵����]� ���������������������U����   SVWQ��4����3   ������Y�M��EP�M��1y��_^[���   ;��0�����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�M�趱��_^[���   ;��д����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�M��M���_^[���   ;��p�����]� ���������������������������U����   SVWQ��4����3   ������Y�M�j �EP�K�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M�j �EP������_^[���   ;�讳����]� �������������������������U����   SVWQ��4����3   ������Y�M�j �EP�]�����_^[���   ;��N�����]� �������������������������U����   SVWQ��4����3   ������Y�M��E����M��B��;������_^[���   ;�������]��������������������U����   SVWQ��4����3   ������Y�M��@QPj �MQ�M��w���_^[���   ;�舲����]� �������������������U����   SVWQ��(����6   ������Y�M��M苉��;Es�M��h����M�v���+E�E�E�;Es�E�E�E��@Q+H;Mw�M��]����} vT�E��HM�M�j �U�R�M��~������t3�EP�M�Y���EP�M��|����M�AP�S������E�P�M������E�_^[���   ;�蕱����]� ����������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��@Q+H;Mw�M��n����} vE�E��HM�M�j �U�R�M��}������t$�EP�MQ�U��BP�M���p���E�P�M��4����E�_^[���   ;�走����]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M�h>  h�V�EP�������EP薝����P�MQ�M�耷��_^[���   ;�������]� ����������������������������������������U����   SVWQ��(����6   ������Y�M��} th*  h�V�EP��������EP�M���o���ȅ�t �EP�M��J����M+�Q�U�R�M��^����n�E��@Q+H;Mw�M�迚���} vL�E��HM�M�j �U�R�M���{������t+�EP�MQ�M������U�BP轤�����E�P�M��~���E�_^[���   ;��������]� ��������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��M�˅��;Es�M�訥���M超��+E�E�E;E�s�E�E�E�;Eu�EE�P�M��6����MQj �M��'����Bj �E�P�M���z���ȅ�t-�E�P�M蝜��EP�M������P蝣�����E�P�M��^~���E�_^[���   ;��߭����]� ����������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E;@Qu�M��Ę��j �EP�M��z���ȅ�t�EP�MQj �M��hm���EP�M��}���E�_^[���   ;��"�����]� ���������������������������������������������U����   SVWQ��4����3   ������Y�M�h�  h�V�EP�������EP������P�MQ�M��9���_^[���   ;�荬����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��} th  h�V�EP�o������EP�M��hl���ȅ�t �EP�M�躓���M+�Q�U�R�M��T����=j �EP�M��x���ȅ�t%�EP�MQ�M�聓��P�^������EP�M��|���E�_^[���   ;�蠫����]� �����������������������������������������������������������U����   SVW��@����0   ������EP�MQ�UR豗����_^[���   ;�������]��������������������������U����   SVW��@����0   ������E�M��_^[��]������������������U����   SVWQ��4����3   ������Y�M��E�P�M��I���P�M�:����E_^[���   ;��t�����]� �������������������������������U����   SVWQ��4����3   ������Y�M��E�P�M��QR�M������E_^[���   ;�������]� ���������������������������������U����   SVWQ��0����4   ������Y�M��E��8 t�M����0�����E�����0�����0���_^[��]��������������������������������U����   SVWQ��4����3   ������Y�M��M��Η��_^[���   ;��4�����]������������������U����   SVWQ��0����4   ������Y�M��E��8 uǅ0����Q��M��	���Ý����0�����0���_^[���   ;�迨����]�����������������������������U����   SVWQ��4����3   ������Y�M��E��M��@+A��0   ��_^[��]�������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��0����4   ������Y�M��E��x8 u�M����0����	�U��0����EP��0���Q�M�賅��_^[���   ;��h�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M�j �M��~w��_^[���   ;�������]��������������������������������U����   SVWQ��4����3   ������Y�M��M�誈���E��HQ�U��BP�M��bt���E��M��Q�P_^[���   ;�肦����]��������������������������������U����   SVWQ��4����3   ������Y�M�j �EP�M��i���_^[���   ;�������]� �������������������������U���P  SVWQ�������T   ������Y�M��E���M��A�E��M��P#Qu��   �E��tj j �,����   �E��M��P#Q��t5j������P訷����Ph(T�������!���h�<������Q�����y�E��M��P#Q��t5j��(���P�b�����PhDT������ۧ��h�<�����Q蝝���3j������P�-�����Ph`T������覧��h�<������Q�h���_^[��P  ;��ؤ����]� �����������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E��E�E��xP u	�E�    �0�M���������u�E�    �E��HPQ�؎������t�E�    jj �M���s���E�_^[���   ;��������]���������������������������������������������������U����   SVWQ��$����7   ������Y�M��EPj0��������,�����,��� t�   �u��,���󥋍,�����$����
ǅ$���    _^[���   ;��G�����]� ����������������������������������U����   SVW��<����1   ������} u�E��<�����MQ�UR�EP�q������<�����<���_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M��t���_^[���   ;��\�����]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M�蜲��_^[���   ;��������]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�MQ�M��;���_^[���   ;�蜡����]� �����������������������U����   SVWQ��4����3   ������Y�M��EP�!�����_^[���   ;��@�����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�������_^[���   ;�������]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�a�����_^[���   ;�耠����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�^������t�����P�EP�M�ph���E���[���P�EP�M�Wh���E_^[���   ;�������]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��E�P�MQ�M��g���E_^[���   ;��y�����]� ��������������������U����   SVWQ��4����3   ������Y�M��_^[��]���������������������U����   SVWQ��4����3   ������Y�M�2�_^[��]���������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M��E�M��U �E��   ��t	�   �D�B��E����U�
�E ����U �
�E�;Mt�E �;Mt�E��U ��	���3�_^[��]� ������������������������������������������������U����   SVWQ��0����4   ������Y�M��E+E9Es�M��0�����U+U��0�����0���_^[��]� ����������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]������������������U����   SVWQ��4����3   ������Y�M��E_^[��]� �����������������U����   SVWQ��4����3   ������Y�M�h
  hR�EP�MQ�n�����h
  hR�EP�b�����E+EP�MQ�UR�<k�����E_^[���   ;��r�����]� ���������������������������������������������U����   SVWQ��4����3   ������Y�M��E�M��U �E��   ��t	�   �D�B��E����U�
�E ����U �
�E�;Mt�E �;Mt�E��U ��	���3�_^[��]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M��E���P�MQ�ي����_^[���   ;��8�����]� �������������������U����   SVWQ��4����3   ������Y�M�h�	  hR�EP�MQ螥�����	�E���E�E;Et�E���P�M�R�J������M��ҋE_^[���   ;�蟚����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��E���P�MQ��l����_^[���   ;��(�����]� �������������������U����   SVWQ��4����3   ������Y�M�h�	  hR�EP�MQ莤�����	�E���E�E;Et�E���P�M�R�\l�����M��ҋE_^[���   ;�菙����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��E�M�3�_^[��]� ��������������������������U����   SVWQ��4����3   ������Y�M��E_^[��]� �����������������U����   SVWQ��4����3   ������Y�M�h�	  hR�EP�MQ�N�����h�	  hR�EP�i^�����E+EP�MQ�UR�g�����E_^[���   ;��R�����]� ���������������������������������������������U����   SVWQ��4����3   ������Y�M��E��H�_^[��]���������������U����   SVWQ��4����3   ������Y�M��E��H�U��B,�	��_^[��]���������������������U����   SVWQ��0����4   ������Y�M��E��x uǅ0���   �
ǅ0���    ��0���_^[��]����������������������������������U����   SVWQ��4����3   ������Y�M��E�P�M��QR�M�͊���E_^[���   ;��֖����]� ���������������������������������U����   SVW��@����0   ��������_^[��]�������������������������U����   SVWQ��4����3   ������Y�M��E��H �U��B0�	��_^[��]���������������������U����   SVW��<����1   ������E�M�;uǅ<���   �
ǅ<���    ��<���_^[��]��������������������U����   SVWQ��0����4   ������Y�M��M����P�M���~������t�M��i��;Euǅ0���   �
ǅ0���    ��0���_^[���   ;��K�����]� ��������������������������������������U����   SVWQ��$����7   ������Y�M��EP��MQ��(���R�E���M��B��;��ה�����z���_^[���   ;��������]� ���������������������������U����   SVWQ��4����3   ������Y�M��E��H;Ms�M�蚋���EP�M���d���E�_^[���   ;��J�����]� �������������������������������������U����   SVWQ������9   ������Y�M��E��H;Ms�M������E��H+M;Mw�EP�M��;d���F�} v@�M��x{��E�E�E��H+M�M��E�+EP�M�MQ�U�R�Sc�����E�P�M���c���E�_^[���   ;��t�����]� �����������������������������������������������U����   SVWQ��0����4   ������Y�M��M���d����tǅ0���   �
ǅ0���    ��0���_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ�� ����8   ������Y���3ŉE��M�E��U�Q���'V����tW�E�P�M������M��͡������t4�E��U�Q����U�����e�����uj j�E��U�Q��������M��c_���E�R��P�l�	�~���XZ_^[�M�3���u�����   ;�跑����]�   t�	����   ��	_Ok ������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��H,�+U�E��H,��E��H�U�E��H�_^[��]� ������������������������������U����   SVW��@����0   ��������_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��E��H4Q�M�ҁ���E_^[���   ;��j�����]� ���������������������U����   SVWQ��4����3   ������Y�M��E��H0Q�M�r����E_^[���   ;��
�����]� ���������������������U����   SVWQ��0����4   ������Y�M��M��a����uǅ0���   �
ǅ0���    ��0���_^[���   ;�蔏����]����������������������������������U����   SVWQ��4����3   ������Y�M��E��H�_^[��]���������������U����   SVWQ��4����3   ������Y�M��EP��q����P�M��i��_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M���M��B��;��*���_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M��M��/U���E��M�H8�E��@<    j �M���z���M��A@�E��x8 uj j�M�蓟���E��t�E�P��Z����_^[���   ;��h�����]� �����������������������������������U����   SVW��@����0   ��������_^[��]�����������������������U����   SVWQ��0����4   ������Y�M��E�M��Q�B�M#�tǅ0���   �
ǅ0���    ��0���_^[��]� ����������������������������������U����   SVW��<����1   ������E���uǅ<���    ��UR��{������<�����<���_^[���   ;��#�����]���������������������������������U����   SVW��@����0   �������g��P�EP�M�Y���E_^[���   ;�輋����]��������������������������U����   SVWQ��4����3   ������Y�M��E�P��h����_^[���   ;��`�����]������������������������������U����   SVWQ��4����3   ������Y�M��E�P豍����_^[���   ;�� �����]������������������������������U����   SVWQ��4����3   ������Y�M����_^[��]��������������������U����   SVWQ��4����3   ������Y�M��UUU_^[��]������������������U����   SVW��@����0   ������M�y���_^[���   ;��)�����]�����������������������U����   SVW��@����0   ������M�t��_^[���   ;��ى����]�����������������������U����   SVWQ������:   ������Y�M���#���P�M���������g���E�}�wǅ���   ��E������������_^[���   ;��O�����]���������������������������������������������U����   SVWQ��(����6   ������Y�M���/���P�M��^����萉��_^[���   ;��ֈ����]��������������������U����   SVWQ��$����7   ������Y�M��EP�g�����E�}� t�E쉅$����
ǅ$����S��$���Q�M�����E_^[���   ;��P�����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��}uh�S�M臏���E���EP�MQ�M��_���E_^[���   ;�过����]� ��������������������������U����   SVWQ��$����7   ������Y�M��EP�&������E�}� t�E쉅$����
ǅ$����S��$���Q�M�����E_^[���   ;��0�����]� �������������������������������������������U����   SVWQ��0����4   ������Y�M��M��Bs����0����M��[����P�EP��0������0����B��;�襆���E_^[���   ;�蒆����]� �����������������������������U����   SVW��<����1   ������} u�E��<�����MQ�UR�EP�4T������<�����<���_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M��xS_^[��]������������������U����   SVWQ��4����3   ������Y�M���S_^[��]������������������U����   SVWQ��4����3   ������Y�M��T_^[��]������������������U����   SVW��8����2   �������|���M9t�U���<����+�|����uǅ8���   �
ǅ8���    ��8�����<�����<���_^[���   ;�跄����]�������������������������������������U����   SVWQ������9   ������Y�M��E��xP u�EP�MQ�UR茁�����E�}� u3��=j�E�P�M�� T���� ���P�M��[���P�g����P�M��/^���� �����E���E�_^[���   ;��������]� ������������������������������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M���M��B��;��j���_^[���   ;��Z�����]� �������������������������������������U����  SVWQ������|   ������Y���3ŉE��M�ǅ����    �z��������EP�����Q��p�����Ѕ�t�EP��s�����3  �W�M��i����t8�M��i�����M��I��;�s"�EP�}�����؋M��Q����E��  ��E�xP u
�z����  �M��zi���E�x@ uL�E�HPQ�UR�p}������P�>D�����ȅ�t�U��������y�������������  �}  �E�   �EP�$}�����E�j j�M���Y���E�P��0���Q�M���w�����ъ�����M��Y���V��D���R�M��w����變��P�E�P�M�Q�U�R�E��HP�M�I@��Y����$�����D�����b����0����b����$������������� ��  �����~������?  �  ��X���P�M��/w�����)����M�+ȉM���X����ab���}� vD�E�HPQ�U�Rj��x���P�M���v��������������P��k����9E�tǅ���   �
ǅ���    �������o�����������t���������x�����a����o�����t�6x���������M���S����������   �E��@E�E�9E�t�E�������M��S���������   �}� v�6�M��{W���� sj j�M��[�����w���������M��|S���������w�h�E�HPQ�U�R��A��������t�M�������w�������������������M��-S���������(�`w���������M��S��������������M���R��R��P���	�+���XZ_^[�M�3��c�����  ;��d����]� �I    ��	����   �	����   �	����   �	����   ��	_Str _Dest _Src _Ch ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��u��_^[���   ;���}����]� ������������������U����   SVW��$����7   �����󫡀�3ŉE�j j�E�P�M�vy���E�E�E�� R��P���	����XZ_^[�M�3��a�����   ;��A}����]Ë�   ��	����   ��	f_buf ��������������������������������������������������U����   SVW������9   ������EP�r�����]��EP�r�����]�EP�}r�����]�Q�E��$Q�E��$Q�E��$�M�	v���E_^[���   ;��h|����]��������������������������������������U���  SVW��������   �����󫡀�3ŉE�h�   ��@����U��jj@j!�M�TI��P��@���������@����H��@����؏���Ѕ�t,j h�U��������W��������P�_�����������c����Q������jOj ������P�h����j jP������P��@����pw��j j������P��@����Zw��������P�������������̍�����P�YU���������%j����������x�����x������l���ǅ`���    ���`�������`�����`���;�l����  ��@���P��L���Q�d������@���P��8���Q�d������@���P��$���Q�d������@���P�����Q�pd�������ċ�����������P������H���ԋ�$������(����J��,����B���̋�8������<����A��@����Q���ċ�L������P����P��T����H������@A��P����������j j�����P��@�����u�������������P�M� N���������I=���������)M����@�����~���ER��P���	�I���XZ_^[�M�3���]����  ;��y����]ÍI 
   ��	@����   Y�	����P   M�	����   A�	����   ?�	����,   :�	L���   3�	8���   0�	$���   -�	���   *�	���   $�	dummy v3 v2 v1 normal info h n_triangles header_info stl_file ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ������?   ������Y�M��M���>������   �M��Z�����M��>��;�s~�/o��������EP�����Q�_e�����Ѕ�u;�M��>���   k���P�|����������EP�����Q�$e�����Ѕ�t�M��s���EP�Bh�����   �   �E��xP t%�n���� ����EP�� ���Q��d�����Ѕ�t	�n���y�w�E��x@ u6�EP��q������/����M��QPR��/���P�H�����ȅ�t�E�:�8�M��=���M���D;�t!�EP�q�����M��AD�M��@���E���n��_^[���   ;��Jv����]� �����������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��em��_^[���   ;��u����]� ������������������U����   SVWQ��4����3   ������Y�M��E��H0�+U�E��H0��E��H �U�E��H �_^[��]� ������������������������������U����   SVWQ��4����3   ������Y�M��E��H �_^[��]���������������U����   SVWQ��4����3   ������Y�M��E����M��B4��;��t��_^[���   ;��t����]��������������������U����   SVWQ������<   ������Y�M��EP�|i����P�M��L���ȅ���   �EP�\i�����M�+A��0   ���E�E��M��P;Qu
j�M��YO���E��HQ�U��BP�M��>��kE�0�M�AP�F<����P�U��BP�����Q�M��I������\���E��H��0�U��J�g�E��M��P;Qu
j�M���N���E��HQ�U��BP�M��=���EP��;����P�M��QR��#���P�M��$I�����d\���E��H��0�U��J_^[���   ;��8s����]� �����������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@8_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U��j�h��d�    PQ��  SVWQ�������B   ������Y���3ŉE�P�E�d�    �e��M�h�  h�W�EP��7�����E�    �E��@    �@    j�E�P�M��P���M��&P��������   �E�    �EP�MQ�UR�E��U�Q���5�����m���E��U��E�HM��PU��E�H�P�E�;Eu�M�;Mt	�E؃��E��jj�E��U�Q���S������	��E�������E�����j �E�P�M��M�J�'����E䉅�����M��i��������R��P�T�	襄��XZ�M�d�    Y_^[�M�3��U����  ;���p����]� ��   \�	����   h�	_Ok ��������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��M�褅����,�����0�����0��� |$	��,��� v�M�����P�t������(�����E����M��B��;���o����(�����(���_^[���   ;��o����]���������������������������������������U����   SVWQ�� ����8   ������Y���3ŉE��M�M��t6���M��D;�u!�}u�E�x@ u�E���M�� �E�M�E�xP tS�M��h������tD�EEu�}t�EP�MQ�UR�E�HPQ�;B������u�E�P�M�QPR�+h������t�4�P�0�Q�M�p>���E�"�M��U���E�P�M�Q�U�BHP�M�cr���ER��P���	�#���XZ_^[�M�3��R�����   ;��\n����]� �I    ��	����   ��	_Fileposition ��������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��4�P�0�Q�M�Y=���E_^[���   ;��m����]� �������������������������������U����   SVWQ������<   ������Y���3ŉE��M�M�ar���E�U�M�@��+E�U�EԉU؋E�xP tb�M��f������tS�E�P�M�QPR�Wb������u<�E�E�tj�E�P�M�Q�U�BPP�@������u�E�P�M�QPR�f������t�4�P�0�Q�M�R<���E�0�M�x1���M�AH�M��S���E�P�M�Q�U�BHP�M�7p���ER��P���	����XZ_^[�M�3��wP�����   ;��0l����]�  �I     �	����   �	_Fileposition ��������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��4�P�0�Q�M�9;���E_^[���   ;��dk����]�  �������������������������������U����   SVWQ��4����3   ������Y�M��M��A�Q_^[��]��������������U����   SVWQ��(����6   ������Y�M��E�P��/���Q�P����P�M�j\���E_^[���   ;��j����]� ������������������������U����   SVWQ��(����6   ������Y�M��E�P��/���Q��V����P�M�A���E_^[���   ;��=j����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�P�M�M���E_^[���   ;���i����]� ������������������������U����   SVWQ��4����3   ������Y�M��E�P�M��P���E_^[���   ;��}i����]� ������������������������U����   SVW��@����0   ������EP�M��4���E_^[���   ;��"i����]��������������������������������U����   SVW��@����0   ������EP�M�)���E_^[���   ;���h����]��������������������������������U����   SVWQ��0����4   ������Y�M��E��xP tF�} u�EEuǅ0���   �
ǅ0���    �MQ��0���R�EP�M��QPR�j������t3���j�E��HPQ�M���7���E�_^[���   ;��h����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ��4����3   ������Y�M��E��H�U��E��H�U��E+E�M��Q,�_^[��]� ��������������������������������U����   SVWQ��4����3   ������Y�M��E��H�U��E��H �U��E+E�M��Q0�_^[��]� ��������������������������������U����   SVWQ��4����3   ������Y�M��} t�EP�M��R8��EP�M��yZ��_^[���   ;��]f����]� ������������������������U����   SVWQ��(����6   ������Y�M��M��{����,�����0�����0��� |$	��,��� v�M��-��P�j������(�����E����M��B��;���e����(�����(���_^[���   ;��e����]���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E���M��B ��;��:e��_^[���   ;��*e����]� �������������������������������������U����   SVWQ��4����3   ������Y�M�3�3�_^[��]�������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��M��@+A��0   ��_^[��]�������������������U����   SVWQ������=   ������Y�M��M��y����������������� |$	�����v�M���M��P�h����������]�M���1���� ����f[����,����� ���P��,���Q�Q�����Ѕ�t�>[���������M��/s����������������������_^[���   ;��Xc����]����������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ������:   ������Y�M��E��xP ti�LZ����P�M���M��B��;��b���� ����*Z����,����� ���Q��,���R�WP��������u�M��QPR�l������}ǅ��������
ǅ���    �����_^[���   ;��b����]��������������������������������������������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]���������������������U����   SVW��@����0   ��������_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��E��@<_^[��]�����������������U����   SVW��@����0   ������E� _^[��]�����������������������U����   SVW��@����0   ������E� _^[��]����������������������U����  SVWQ�� ����x   ������Y���3ŉE��M�M��'����t.�M��'�����M��cB��;�s�M��=u��P�e�����  ��E�xP u
��W���  �M��6G���E�x@ uM�E� �E�HPQ�U�R��8��������t�M�Q�d������ �����W���� ����� ����L  �G  �M��	p���E�HPQ�4 �����E��}��u�PW����(����M��3����(����	  �E�Pj�M���:���E�P�M�Q�U�R�E�P��@���Q�M��[U�����Uh�����M��6���V��T���R�M��8U�����2h��P�E��HP�M�I@�X����4�����T����Y@����@����N@����4����� ����� ��� �A  �� ���~�� �����   �&  �E�9E���   ��h���P�M��T�����g�����M���5���+u��u���h�����?���}� ~$�E����E��M�QPR�E�E��Q��N�����֍E�P�%c������|����M��1����|�����   �1������P�M��/T�����)g���M�+�Qj �M��	O���������Y?���~�M��J5����s�oj������P�M���S������f��Pj�M�Q�C/�����������?���E�P�b�����������M��1���������(�QU���������M��1���������������M���0��R��P��
�q��XZ_^[�M�3��A�����  ;��U]����]Ë�   �
����   (
����   #
����   
����   
����   
_Src _Dest _Ch _Str _Ch ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ������:   ������Y�M��E����M��B��;���[���� ����iS����,����� ���Q��,���R�I��������t�AS���������M��xp��P�F`��������������_^[���   ;��^[����]��������������������������������������������U����   SVWQ������:   ������Y���3ŉE��M�M��$"����t+�M��"�����M���<��;�s�M��"��P�_�����d�b�E���M�B��;��Z���E��[R��������M�Q�����R�H��������t�E�����E�P�M��M�B��;��lZ���E�R��P��
�n��XZ_^[�M�3��>�����   ;��>Z����]ÍI    �
����   �
_Meta ������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��UQ��_^[���   ;��Y����]���������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M���M��B ��;��6Y��_^[���   ;��&Y����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ������9   ������Y�M��� ���P�M��PA��P��<�����E썍 ����)���EP�M��e��_^[���   ;��X����]� ������������������������������������U����   SVWQ��4����3   ������Y�M����EP�M���M��B ��;��W��_^[���   ;��W����]� ����������������������������U���  SVWQ�������B   ������Y���3ŉE��M�fW�fEȃ} �"  
�} �  �M��l���E؉U܃}� |}�}� vu�E;E�|�M;M�s�E�E؋M�M܋E�P�M����P�MQ�L�����E�E�E�E�E؋M�M܉EȉM̋E+E؋MM܉E�M�E�P�M��{���   �E���M�B��;��V���E��2N���������M�Q������R�bD��������t�E�>�E�P�Q�����M��U���U�Eȃ��M̃� �EȉM̋E���M�� �E�M������EȋU�R��P�<

�i��XZ_^[�M�3��3:����  ;���U����]� �I    D

����   P

_Meta ��������������������������������������������������������������������������������������������������������������������������U���  SVWQ�������A   ������Y�M�fW�fE؃} �$  
�} �  �M��B���E�U�}� |}�}� vu�E;E�|�M;M�s�E�E�M�M�E�P�MQ�M��;��P�YJ�����E�E�E�E�E�M�M�E؉M܋E+E�MM�E�M�E�P�M��a8���   �EP�<Y������P�M���M��B��;��YT���� �����K��������� ���Q�����R�)B��������t�4�-�E���E�E؃��M܃� �E؉M܋E���M�� �E�M������E؋U�_^[��  ;���S����]� ����������������������������������������������������������������������������������������������������������U����   SVW��@����0   ��������E�$���E�$�[����_^[���   ;��S����]�����������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��NR����E�P�MQ����B�H�у�;��,R���E�_^[���   ;��R����]� ������������������������������������U����   SVWQ��4����3   ������Y�M��M���C��_^[���   ;��Q����]������������������U����   SVWQ��0����4   ������Y�M��EP�M��Pb����uǅ0���   �
ǅ0���    ��0���_^[���   ;��@Q����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M��P���E��t�E�P�d�����E�_^[���   ;���P����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bx��;��nP��_^[���   ;��^P����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��PH��;���O��_^[���   ;���O����]� �������������������������������������U����   SVWQ������:   ������Y�M��E��x t�   �E��8 t)��E��Q����B<�H�у�;��fO���E��     �E��x tS�E��x t@�E��H��,�����,����� ����� ��� tj�� �����E��������
ǅ���    �E��@    _^[���   ;���N����]���������������������������������������������������������������U����   SVW��@����0   ���������@��_^[���   ;��wN����]���������������������U���x  SVW�������^   ������EP����q3��P�M��*��j h�^�������F*��j �E�P������Q�M��'����uǅ����   �
ǅ����    ��������������������5����������t�M�S���M���5���E�  j�E�P�M��O��j�j��EP�M�Q�M��L��j h�^�������)��j �E�P������Q�M��o&����uǅ����   �
ǅ����    �������������������M5����������t�M��R���M��25���E�p  j�E�P�M����j�j��EP�M�Q�M���K��j h�^�������)��j �E�P������Q�M���%����uǅ����   �
ǅ����    �������������������4����������t�M�HR���M��4���E��   j�E�P�M����j�j��EP�M�Q�M��OK��j h�^������o(��j �E�P�����Q�M��5%����uǅ����   �
ǅ����    ������������������4����������t�M�Q���M���3���E�9j�E�P�M��{��j�j��EP�M�Q�M��J���E�P�M�:(���M��3���ER��P��
�>_��XZ_^[��x  ;��K����]Ë�   �
����   �
����   �
str pos ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���T  SVW�������U   ������EP����/��P�M���&��j h�^�������v&��j �E�P������Q�M��<#����uǅ����   �
ǅ����    �������������������2����������t�M�O���M���1���E�p  j�E�P�M����j�j��EP�M�Q�M��H��j h�^��������%��j �E�P������Q�M��"����uǅ����   �
ǅ����    �������������������}1����������t�M�O���M��b1���E��   j�E�P�M�����j�j��EP�M�Q�M��H��j h�^������<%��j �E�P�����Q�M��"����uǅ����   �
ǅ����    �������������������0����������t�M�xN���M���0���E�9j�E�P�M��H��j�j��EP�M�Q�M��G���E�P�M�%���M��0���ER��P��
�\��XZ_^[��T  ;��NH����]ÍI    �
����   �
����   �
str pos ����������������������������������������������������������������������������������������������������������������������������������������������������������������U���0  SVW�������L   ������EP����,��P�M���#��j h�^�������f#��j �E�P������Q�M��, ����uǅ����   �
ǅ����    �������������������
/����������t�M�L���M���.���E��   j�E�P�M��o��j�j��EP�M�Q�M��E��j h�^�������"��j �E�P�����Q�M������uǅ����   �
ǅ����    ������������������m.����������t�M�L���M��R.���E�9j�E�P�M�����j�j��EP�M�Q�M��E���E�P�M�"���M��.���ER��P�H
�Y��XZ_^[��0  ;���E����]�   P
����   l
����   h
str pos ��������������������������������������������������������������������������������������������������������������������������������U���  SVW�������C   ������EP����A*��P�M��!��j h�^������!��j �E�P�����Q�M�������uǅ����   �
ǅ����    ������������������,����������t�M�RJ���M��,���E�9j�E�P�M��"��j�j��EP�M�Q�M��\C���E�P�M�� ���M��d,���ER��P��
��W��XZ_^[��  ;��(D����]Ð   
����    
����   
str pos ��������������������������������������������������������������������������������������������U����   SVW��@����0   ������EP����(��_^[���   ;��cC����]�����������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BT�Ѓ�;���B��_^[���   ;��B����]�������������������������U����   SVW��@����0   �������EP����Q<�B�Ѓ�;��cB��_^[���   ;��SB����]���������������������������������U����   SVWQ������9   ������Y�M���EP�MQ�� ���R����P�M����   ��;���A��P�M�e���� �����)���E_^[���   ;��A����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BH�Ѓ�;��KA��_^[���   ;��;A����]�������������������������U����   SVWQ��$����7   ������Y�M��E��x ufh�^����Ph��j��������,�����,��� t�MQ��,����@J����$����
ǅ$���    �U���$����B�E��x u3���E��x t&�E��8 tǅ$���   �
ǅ$���    ��$����P��EP����Q<��Ѓ�;��A@���M���E��@   �E��8 tǅ$���   �
ǅ$���    ��$���_^[���   ;���?����]� �������������������������������������������������������������������������U����   SVWQ������?   ������Y�M������P�N+����P�M��H/��������������������_^[���   ;��M?����]���������������������������U����   SVWQ��0����4   ������Y�M��E��@   ����H<��Q��;���>���M���E��8 tǅ0���   �
ǅ0���    ��0���_^[���   ;��>����]���������������������������������U����   SVWQ��4����3   ������Y�M��E��8 u����H��#��EP�M��R����H<�Q�҃�;��5>��_^[���   ;��%>����]� ��������������������������������U����   SVW��<����1   ������} t�E��<�������������<�����<���Q�UR�EP�5����_^[���   ;��=����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E��x t�   �4�E��x u3��'��E��HQ�U��P����Q<�B�Ѓ�;��=��_^[���   ;���<����]��������������������������������������U����   SVW������:   ������} u3��   �EP�M�����E�    �E�    �E�P�M�Q�M��<����tT�}�t�}�u"�EP�M��-��P��Q������t�   �*�$�}�u�EP�M��%�����N����t�   ��3�R��P�$$
�O��XZ_^[���   ;���;����]�   ,$
����   W$
����   T$
����   P$
dat id browse ����������������������������������������������������������������������������������U���p  SVW�������\   ������ǅ����    j h�^�������c��P��M�����E��������6#���}� u3���   �E�    �E�P�M�����E�P�M�Q�M��*;������   �}���   �M�����E��}� tF�EP�������@��������Pj������Q�M��F������������L����tǅ����   �
ǅ����    ��������������������t��������������j"����������t��������������M"����������t�EԉE�������E�R��P�,&
�M��XZ_^[��p  ;���9����]Ë�   4&
����   c&
����   _&
����   X&
browse dat id ��������������������������������������������������������������������������������������������������������������������������U���d  SVW�������Y   ������ǅ����    �} u6j h�^�������-��P�K�����E������� !���} u3��$  �E�    �EP�M��� ���E�P�M�Q�M���8������   �}���   �M��m ���Eă}� tF�EP�������I>��������Pj������Q�M��������������J����tǅ����   �
ǅ����    ��������������������t��������������4 ����������t�������������� ����������t�E��E��2�+�}�u%�}� t�EP�M�� �����1J����t�E��E��������E�R��P��(
�SK��XZ_^[��d  ;��7����]ÍI    �(
����   �(
����   �(
����   �(
browse dat id ��������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �����󫡸��H<��Q��;��6��_^[���   ;��6����]�������������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;��6���j�EP�
  ��_^[���   ;���5����]���������������������������������������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;��E5���j�EP��	  ��_^[���   ;��%5����]���������������������������������������������������U����   SVW��<����1   ������=�� tI�}sǅ<���   �	�E��<�����MQ�UR��<���P����Q���   �Ѓ�;��4���j�EP�	  ��_^[���   ;��a4����]�����������������������������������������������U����   SVW��<����1   ������=�� ��   �} tK�}sǅ<���   �	�E��<�����MQ�UR��<���P����Q���   �Ѓ�;��3���[�I�}sǅ<���   �	�E��<�����MQ�UR��<���P����Q���  �Ѓ�;��l3����EP�MQ��  ��_^[���   ;��J3����]������������������������������������������������������������������������U����   SVW��4����3   ������} tN�E�E��=� t"�   k���U�<
�u�E��P�@=�������E�P����Q��Ѓ�;��2��_^[���   ;��}2����]�������������������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��2��_^[���   ;��2����]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��1��_^[���   ;��1����]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��41��_^[���   ;��$1����]����������������������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;��0���j�EP�)  ��_^[���   ;��u0����]���������������������������������������������������U����   SVW��<����1   ������=�� tE�}sǅ<���   �	�E��<�����j j ��<���Q����B���   �у�;���/���j�EP�i  ��_^[���   ;��/����]���������������������������������������������������U����   SVW��0����4   ������} w�E   �=�� t0��EP�MQ�UR����H���   �҃�;��#/����0����j�EP�  ����0�����0����M��E���th _����
P�m@�����E�_^[���   ;���.����]�����������������������������������������������������������U����   SVW��0����4   ������} w�E   �=�� to�} t0��EP�MQ�UR����H���   �҃�;��-.����0����.��EP�MQ�UR����H���  �҃�;���-����0�����0����E��j�EP�  ���E��E���th _����P�J?�����E�_^[���   ;��-����]������������������������������������������������������������������������U����   SVW��4����3   ������} tN�E�E��=� t"�   k���U�<
�u�E��P�7�������E�P����Q��Ѓ�;���,��_^[���   ;���,����]�������������������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��t,��_^[���   ;��d,����]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��,��_^[���   ;���+����]����������������������������������U����   SVW��@����0   �������EP����Q��Ѓ�;��+��_^[���   ;��+����]����������������������������������U����   SVW��4����3   ������}s�E   �E��P�������E��}� u3��:�} t�E��Pj �M�Q������E�� �����E����E���   �E�_^[���   ;���*����]��������������������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��\*��_^[���   ;��L*����]��������������������������U����   SVW��@����0   �������EP�MQ����B��  �у�;���)��_^[���   ;���)����]��������������������������U����   SVW��@����0   �����󫡸��H��   ��;��)��_^[���   ;��x)����]����������������������U����   SVW��@����0   ������} t�   k���U�<
�u�   �3�_^[��]����������������������������U����   SVW��@����0   ������} t!��EP����Q��@  �Ѓ�;��(��_^[���   ;��(����]������������������������U����   SVW��@����0   �������hﾭޡ���H��@  �҃�;��P(��_^[���   ;��@(����]������������������������������U����   SVW��@����0   ������E�8 t��E�Q����B��у�;���'���E�     _^[���   ;���'����]�������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��j �EP�M�Q������   �H�у�;��B'���E�_^[���   ;��/'����]� ������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   ��Ѓ�;��&��_^[���   ;��&����]��������������������������U����   SVWQ��4����3   ������Y�M��E���P�)����_^[���   ;��M&����]���������������������������U����   SVW��(����6   ������EP�M�����EP�M��82���E�P�M�z���M������ER��P�d:
�~9��XZ_^[���   ;���%����]Ë�   l:
����   x:
s ��������������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��@%��_^[���   ;��0%����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B�Ѓ�;���$��_^[���   ;��$����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B�Ѓ�;��B$��_^[���   ;��2$����]� �����������������������������U����   SVW��@����0   �����󫡸��H0�􋑤   ��;���#��_^[���   ;���#����]����������������������U����   SVW��@����0   �����󫡸��H8����;��|#��_^[���   ;��l#����]��������������������������U����   SVW��@����0   �����󫡸��H8��Q<��;��#��_^[���   ;��#����]�������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q���  �Ѓ�;��"��_^[���   ;��"����]����������������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ����B��  �у� ;��"��_^[���   ;��"����]����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B,�Ѓ�;��!��_^[���   ;��!����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q8�B4�Ѓ�;��!��_^[���   ;��!����]� �����������������������������U����   SVW������=   �������2����u�\h���M������EPh���M��j���EPh���M��Y��j �E�PhicMC�����Q�%%����������5����M�����R��P��?
��3��XZ_^[���   ;��9 ����]Ë�   �?
����    @
msg ������������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��l  �҃�;����_^[���   ;������]�����������������������U����   SVW��@����0   �������EP����Q��\  �Ѓ�;��0��_^[���   ;�� ����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q0���   �Ѓ�;����_^[���   ;������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B8�HD�у�;��J��_^[���   ;��:����]� �������������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ����B��$  �у�;��\��_^[���   ;��L����]��������������������������U����   SVW��@����0   �������EP�MQ����B�Hx�у�;�����_^[���   ;�������]�����������������������������U����   SVW��@����0   �����󫡸��H���  ��;����_^[���   ;��x����]����������������������U����   SVW��@����0   �������EP���E�$���E�$�MQ����B���   �у�;����_^[���   ;�������]��������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E�P����Q8�B�Ѓ�;��v��_^[���   ;��f����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H8�Q�҃�;�����_^[���   ;�������]� ��������������������������������������U����   SVW��@����0   �������EP����Q��D  �Ѓ�;��p��_^[���   ;��`����]������������������������������U����   SVW��@����0   �������EP����Q��H  �Ѓ�;�� ��_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;����_^[���   ;��y����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;����_^[���   ;��	����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;����_^[���   ;������]�����������������������U����   SVW��@����0   �����󫡸��H�􋑄   ��;��H��_^[���   ;��8����]����������������������U����   SVW��(����6   �������j �EP�MQ�UR�EP��,���Q����B��t  �у�;�����P�M�O�����,���������E_^[���   ;������]����������������������������������U����   SVW��@����0   �������EP������   ���   �Ѓ�;��=��_^[���   ;��-����]���������������������������U����   SVW��@����0   �������E�Q����B0���   �у�;������E�     _^[���   ;������]�����������������������������������U����   SVW��@����0   �������E�Q����B8�H�у�;��Q���E�     _^[���   ;��8����]��������������������������������������U����   SVW��@����0   �������E�Q����B8�H@�у�;������E�     _^[���   ;������]��������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��x  �Ѓ�;��D��_^[���   ;��4����]����������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;�����_^[���   ;������]��������������������������U����   SVW��@����0   �������EP�MQ����B�HP�у�;��_��_^[���   ;��O����]�����������������������������U����   SVW��@����0   �������EP����Q��,  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW������<   ������EPj h�_���������P�M�Q�����������������E�P����Q�B�Ѓ�;��U���M��e���R��P��L
��&��XZ_^[���   ;��,����]Ð    M
����   M
s ��������������������������������������������������U����   SVW��4����3   ������j �M����E��}� t�E�P������E�P������R��P��M
�2&��XZ_^[���   ;��u����]Ë�   �M
����   �M
c ������������������������������������������U����  SVW��(����6  �����󫡀�3ŉE��E�E�E�P�MQh   ������R�����������Ph�_����Q��4  �Ѓ�;�����E�    R��P��N
�Q%��XZ_^[�M�3���������  ;������]ÍI    �N
����   �N
t ��������������������������������������������������������������U����   SVW��@����0   �������EP����Q��8  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �����󫡸��H��QH��;����_^[���   ;��{����]�������������������������U����   SVW��@����0   �����󫡸��H��QD��;��+��_^[���   ;������]�������������������������U����   SVW��@����0   �����󫡸��H��Q<��;�����_^[���   ;������]�������������������������U����   SVW������9   ������EP��MQ�� ���R����H��t  �҃�;��V�����M ���� ��������E_^[���   ;��1����]�������������������������������U����   SVW��(����6   �������,���P����Q��  �Ѓ�;�����P�M�Q�����,���������E_^[���   ;������]������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H�QL�҃�;��<��_^[���   ;��,����]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q���  �Ѓ�;�����_^[���   ;������]����������������������������������U����   SVW��(����6   ������M��,����E�P����Q�B8�Ѓ�;��K���E�P�M������M��O����ER��P�S
�� ��XZ_^[���   ;������]�   S
����   $S
str ����������������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;����_^[���   ;������]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;����_^[���   ;��	����]�����������������������U����   SVW��(����6   �������,���P����Q��  �Ѓ�;����P�M�1�����,��������E_^[���   ;������]������������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����Q���  �Ѓ�;����_^[���   ;���
����]��������������������������������������U����   SVW��@����0   ������E��P��P�M��@Q�U��0R�E�� P�M��Q�UR�EP����Q���   �Ѓ�;��i
��_^[���   ;��Y
����]���������������������������������������U����   SVW��@����0   �����󫡸��H���  ��;���	��_^[���   ;���	����]����������������������U����   SVW��@����0   �����󫡸��H�􋑼   ��;��	��_^[���   ;��	����]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B���  �у�;�� 	��_^[���   ;��	����]������������������������������U����   SVW��@����0   �������EP����Q��L  �Ѓ�;����_^[���   ;������]������������������������������U����   SVW��@����0   ������E�8 t#��E�Q����B��D  �у�;��6���E�     _^[���   ;������]���������������������������U����   SVW��@����0   �������EP�MQ�UR����H��X  �҃�;����_^[���   ;������]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H��\  �҃�;��I��_^[���   ;��9����]�����������������������U����   SVW��@����0   �������EP����Q��H  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR����H���  �҃�;��]��_^[���   ;��M����]���������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ�UR����H���  �҃�;�����_^[���   ;�������]���������������������������U����   SVW��@����0   �������EP�MQ�UR����H��P  �҃�;��i��_^[���   ;��Y����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H��T  �҃�;�����_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H��@  �҃�;����_^[���   ;��y����]�����������������������U����   SVW��@����0   �����󫡸��H���  ��;��(��_^[���   ;������]����������������������U����   SVW��@����0   �����󫡸��H��p  ��;�����_^[���   ;������]����������������������U����   SVW��@����0   �������EP����Q��<  �Ѓ�;��`��_^[���   ;��P����]������������������������������U����   SVW��@����0   �������EP�MQ����B�H@�у�;�����_^[���   ;�������]�����������������������������U����   SVW��@����0   �������EP�MQ����B��  �у�;��|��_^[���   ;��l����]��������������������������U����   SVW��@����0   �������EP����Q�B�Ѓ�;����_^[���   ;������]���������������������������������U����   SVW��@����0   �������EP����Q��\  �Ѓ�;����_^[���   ;������]������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��0��_^[���   ;�� ����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQh�2  ����B���   �у�;�� ��_^[���   ;�� ����]�����������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���   �҃�;��) ��_^[���   ;�� ����]�����������������������U����   SVW��@����0   �������EP�MQ����B���   �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;��P���_^[���   ;��@�����]������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;��p���_^[���   ;��`�����]������������������������������U����   SVW��@����0   �������EP�MQ����B���   �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP�MQ����B��|  �у�;�����_^[���   ;��|�����]��������������������������U����   SVW��@����0   �������EP����Q�B,�Ѓ�;��#���_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP����Q��T  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��<���_^[���   ;��,�����]��������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��  �Ѓ�;������_^[���   ;�������]����������������������������������U����   SVW��@����0   �����󫡸��H��P  ��;��X���_^[���   ;��H�����]����������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��d  �Ѓ�;������_^[���   ;��������]����������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVW��@����0   �������EP����Q��,  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �����󫡸��H��<  ��;�����_^[���   ;��x�����]����������������������U����   SVW��@����0   �����󫡸��H��0  ��;��(���_^[���   ;�������]����������������������U����   SVW������=   �������R�����u�M�����E�^h����M�������EPh����M�����j �E�PhicMC�����Q�K��������g���P�M����������K����M�������ER��P��g
�	��XZ_^[���   ;��L�����]Ð   �g
����   �g
msg ����������������������������������������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW������=   �������������u�M�����E�^h!���M��l����EPh!���M������j �E�PhicMC�����Q��������������P�M���������������M��@����ER��P�Xi
�
��XZ_^[���   ;��������]Ð   `i
����   li
msg ����������������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��`  �҃�;��)���_^[���   ;�������]�����������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P����Q���   �Ѓ�;�������u3���E�R��P��j
�@	��XZ_^[���   ;�������]�   �j
����   �j
����   �j
����   �j
data sub_id main_id ������������������������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW������9   ������M��v�����E�P�MQ����B�H|�у�;��W����E�P�M������M�蟻���ER��P�l
����XZ_^[���   ;�������]�   l
����   l
fn �����������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �B8�Ѓ�;�����_^[���   ;��{�����]�������������������������U����   SVW������=   ������j hLGOg������]���PhicMC�E�P�������������b����M��ٺ����u�M�P����M�������E��M�踺��P�M������M������ER��P�pm
�q��XZ_^[���   ;�������]Ð   xm
����   �m
dat ��������������������������������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P����Q���   �Ѓ�;�������u3���E�R��P�@n
���XZ_^[���   ;��������]�   Hn
����   xn
����   qn
����   ln
data sub_id main_id ������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q0���   �Ѓ�;��+���_^[���   ;�������]�������������������������U����   SVW��(����6   �������EP��,���Q����B���  �у�;�����P�M�=�����,��������E_^[���   ;�������]��������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��0���_^[���   ;�� �����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B8�H �у�;�����_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B0���   �у�;��+���_^[���   ;�������]� ��������������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��$����7   �������EP��(���Q����B���  �у�;��9���P�M�-�����(����u����E_^[���   ;�������]��������������������������������U����   SVW��@����0   �����󫡸��H�􋑄  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������EP����Q��(  �Ѓ�;��P���_^[���   ;��@�����]������������������������������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P����Q���   �Ѓ�;��������u3���E�R��P��s
�` ��XZ_^[���   ;�������]�   �s
����   �s
����   �s
����   �s
data sub_id main_id ������������������������������������������������U����   SVW��@����0   �������EP�MQ����B��l  �у�;������_^[���   ;��������]��������������������������U����   SVW��(����6   �������EP��,���Q����B���  �у�;��y���P�M�������,����}����E_^[���   ;��R�����]��������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������EP�MQ����B��l  �у�;��|���_^[���   ;��l�����]��������������������������U����   SVW�� ����8   �������EP��$���Q����B���   �у�;��	����U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��������]�����������������������������������������������U����   SVW��$����7   ������M��˫����E�P����Q���   �Ѓ�;��X����E�P�M�I����M�蔭���ER��P�w
�����XZ_^[���   ;�� �����]Ð   w
����   w
bc �����������������������������������������������������U����   SVW��@����0   �����󫡸��H��`  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������EP����Q��   �Ѓ�;��0���_^[���   ;�� �����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H8�Q$�҃�;�����_^[���   ;�������]� ��������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��)���_^[���   ;�������]�����������������������U���   SVW�� ����@   �������R�����u3��^hs���M�������EPhs���M�����j �E�PhicMC�����Q�T��������Z��������������W����M��̪�������R��P��y
����XZ_^[��   ;��U�����]Ë�   �y
����   �y
msg ��������������������������������������������������������U���   SVW�� ����@   �������R�����u3��^h#���M�������EPh#���M�����j �E�PhicMC�����Q�T��������Z��������������W����M��̩�������R��P��z
����XZ_^[��   ;��U�����]Ë�   �z
����   �z
msg ��������������������������������������������������������U����   SVW��@����0   �������EP�MQ����B��h  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��L���_^[���   ;��<�����]��������������������������U����   SVW��@����0   �������E$P�M Q�UR�EP�MQ�UR�EP�MQ����B���  �у� ;������_^[���   ;�������]����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H8�Q(�҃�;��G���_^[���   ;��7�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H8�Q0�҃�;������_^[���   ;�������]� ����������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���   �҃�;��I���_^[���   ;��9�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;������_^[���   ;��������]�����������������������U����   SVWQ��4����3   ������Y�M���E�P����Q8�B�Ѓ�;��n���_^[���   ;��^�����]����������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�� ���_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H8�Q�҃�;�����_^[���   ;��w�����]� ����������������������������������U����   SVW��@����0   �������EP����Q��8  �Ѓ�;�����_^[���   ;�� �����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B8�H8�у�;�����_^[���   ;�������]� �������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;�����_^[���   ;��	�����]�����������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��(����6   �������EP�MQ�UR��,���P����Q��X  �Ѓ�;��1���P�M�������,��������E_^[���   ;��
�����]����������������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����Q��h  �Ѓ�;�����_^[���   ;��x�����]��������������������������������������U����   SVW��@����0   �����󫡸��H��d  ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �������EP�MQ����B��@  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ����B���   �у�;��<���_^[���   ;��,�����]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��P4��;������_^[���   ;�������]� �������������������������������������U����   SVW��@����0   �������EP����Q�BT�Ѓ�;��S���_^[���   ;��C�����]���������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;������_^[���   ;��������]��������������������������U����   SVW��@����0   �������EP����Q��  �Ѓ�;��p���_^[���   ;��`�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��  �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP����Q�BX�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP����Q�B\�Ѓ�;��#���_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H�Qt�҃�;��<���_^[���   ;��,�����]��������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M舨��P�U�R����H0���   �҃�(;�����_^[���   ;�������]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�d���P�U�R����H0���   �҃�(;������_^[���   ;��������]�$ ����������������������������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P����Q0���   �Ѓ�(;��G���_^[���   ;��7�����]�$ ����������������������������������U����   SVW��@����0   �������E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR����H���  �҃�$;�����_^[���   ;�������]�������������������������������U����   SVW��@����0   �����󫡸��H��Qd��;��K���_^[���   ;��;�����]�������������������������U����   SVW��@����0   �������EP����Q�Bl�Ѓ�;������_^[���   ;��������]���������������������������������U����   SVW��@����0   �����󫡸��H��Qh��;��{���_^[���   ;��k�����]�������������������������U����   SVW��@����0   �������EP����Q�Bp�Ѓ�;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �����󫡸��H��Q`��;�����_^[���   ;�������]�������������������������U����   SVW��(����6   �������EP�MQ�UR�EP��,���Q����B���  �у�;��-���P�M�������,��������E_^[���   ;�������]������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H0���   �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B0���   �у�;�����_^[���   ;��������]� ��������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���   �҃�;�����_^[���   ;��y�����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;�����_^[���   ;��	�����]�����������������������U����   SVW��4����3   ������} 3��^�EP�MQ�UR�EP�������E��}� |�E��9E�|/�}� }hP_����P�������EE�@� �E���E��E�_^[���   ;��Y�����]���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M��Bh��;������_^[���   ;��������]� ����������������������������������U����   SVWQ������9   ������Y�M���EP����Q�M��Bd��;��n����E�}� u3��s��h�_����P�M��Q����B���   �у�;��/����E��}� u3��4��EP�M��Q�U�R����P�M��Bh��;�������E�E��  �E�_^[���   ;��������]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��Bx��;��`���_^[���   ;��P�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��B��;������_^[���   ;��������]� ����������������������U����   SVW��(����6   �������EP��,���Q����B�H(�у�;��|���P�M� �����,���耵���E_^[���   ;��U�����]�����������������������������������U���  SVW�������`   ������} ��   	�}   @v~j h`����������Pj0j jj �E�U��+�����菵���^`���$������P�9�����P�MQ�>�����������讴��������裴���E�_  �  �} ��   	�}   v{j h`������腨��Pj0j jj �E�U�
������������^`���$������P覷����P�MQ諯�������������������������E��   �~�} |x	�}   vmj h`�����������Pj0j jj �U�M�y����^`���$������P�#�����P�MQ�(�����������蘳��������荳���E�Lj h`�����茧��P�EP��,���Q������P�UR�ڮ������,����J���������?����E_^[�Ā  ;�������]��������������������������������������������������������������������������������������������������������������������������������������������������U���  SVW�������E   �����󫡀�3ŉE��E�E��E�    �E��D�0�Mԃ��MԋE��D�x�Mԃ��M��E�   �	�Eȃ��Eȃ}� |I�E�M������E��E���
}�E���0�MԈD��Uԃ��U���E���7�MԈD��Uԃ��U�먋Eԉ�����������s�������������D� j �E�P�M�å���ER��P���
�.���XZ_^[�M�3�训����  ;��g�����]�   Ė
����   Ж
hexstring ��������������������������������������������������������������������������������������U����   SVW��(����6   ��������E P�MQ�UR�EP���E�$��,���Q����B�H$�у�;�����P�M������,���薰���E_^[���   ;��k�����]�����������������������������������������U����   SVW��(����6   ������j h�  h���,���P�M�������������,���������_^[���   ;��������]�����������������������������U����   SVW��@����0   ������j h�  h��M������_^[���   ;��x�����]����������������������U����   SVW��(����6   ������j h�  h���,���P�M�$�����������,����,�����_^[���   ;��������]�����������������������������U����   SVW��@����0   ������j h�  h��M������_^[���   ;�������]����������������������U����   SVW��@����0   ������h� �M�������tj h�  h��M�T������0����h�_h��k�������_^[���   ;�������]������������������������������������������U����   SVWQ��4����3   ������Y�M��E�� (`�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E�� (`_^[��]��������������U����   SVWQ��4����3   ������Y�M��M��׷���E��t�E�P��������E�_^[���   ;��������]� ������������������������U����   SVW��@����0   �������EP�MQ����B��x  �у�;�����_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ����B��p  �у�;��,���_^[���   ;�������]��������������������������U����   SVWQ������=   ������Y�M��E��E�}� tM�E쉅 ����� ������������� t%��j��������������;�����������
ǅ���    �E�    _^[���   ;��l�����]������������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ����B��  �у�;�����_^[���   ;��|�����]��������������������������U����   SVWQ������<   ������Y�M������P����Q�M���   ��;�����P�M����������`����E_^[���   ;��������]� ��������������������������������������������U����   SVW��@����0   �����󫡸��H��  ��;�����_^[���   ;��x�����]����������������������U����   SVWQ��4����3   ������Y�M�����P��M���$  ��;�� ���_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M�����P��M���(  ��;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �����󫡸��H��d  ��;��H���_^[���   ;��8�����]����������������������U����   SVWQ��4����3   ������Y�M�����P��M���  ��;�����_^[���   ;��п����]������������������������������U����   SVW��@����0   �������EP����Q���  �Ѓ�;��p���_^[���   ;��`�����]������������������������������U����   SVW��@����0   �������EP����Q��|  �Ѓ�;�� ���_^[���   ;�������]������������������������������U����   SVW��@����0   �������EP�MQ����B��t  �у�;�茾��_^[���   ;��|�����]��������������������������U����   SVWQ��4����3   ������Y�M��M��������E�P����Q$�BD�Ѓ�;�������E�P�MQ����B$�HL�у�;�������E�_^[���   ;�������]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��G�����E�P����Q$�BD�Ѓ�;��f�����EP�M�Q����B$�H�у�;��D����E�_^[���   ;��1�����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M�������E�P����Q$�BD�Ѓ�;�趼����EP�M�Q����B$�Hd�у�;�蔼���E�_^[���   ;�聼����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��M��������E�P����Q$�BD�Ѓ�;������E�_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�BH�Ѓ�;�莻���M�螣��_^[���   ;��v�����]������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B$�HL�у�;��
����E�_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B�H�у�;�芺���E�_^[���   ;��w�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H<�у�;��
���_^[���   ;��������]� �������������������������������������U����   SVWQ��0����4   ������Y�M���EP�M�Q����B$�H<�у�;�芹����uǅ0���   �
ǅ0���    ��0���_^[���   ;��Z�����]� �������������������������������������U����   SVW������9   ������EP�M�������EP�M�Q����B$�H@�у�;������E�P�M�_����M��+����ER��P�x�
�h���XZ_^[���   ;�諸����]�   ��
����   ��
fn �������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H@�у�;������E�_^[���   ;�������]� ����������������������������������U����   SVW��@����0   �����󫡸��H(��Q��;�諷��_^[���   ;�蛷����]�������������������������U����   SVW��@����0   �����󫡸��H(����;��L���_^[���   ;��<�����]��������������������������U����   SVW��@����0   �������j j ����H,��҃�;�����_^[���   ;��ն����]�����������������������������������U����   SVW��@����0   �����󫡸��H,��Q,��;��{���_^[���   ;��k�����]�������������������������U����   SVW��@����0   �����󫡸��H���   ��;�����_^[���   ;�������]����������������������U����   SVW��@����0   �����󫡸��H$��QX��;�軵��_^[���   ;�諵����]�������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B(�H�у�;��C���_^[���   ;��3�����]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H0�у�;��ʴ��_^[���   ;�躴����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�B(�Ѓ�;��N���_^[���   ;��>�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�Bh�Ѓ�;��޳��_^[���   ;��γ����]����������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B��;��s���_^[���   ;��c�����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P��M��B��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q$�B�Ѓ�;�莲��_^[���   ;��~�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�HL�у�;�����_^[���   ;��
�����]� �������������������������������������U����   SVW��(����6   �������EP�MQ��,���R����H���  �҃�;�薱��P�M������,���蚙���E_^[���   ;��o�����]���������������������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;������_^[���   ;�������]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;�艰��_^[���   ;��y�����]�����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q$�M��B��;�����_^[���   ;�������]� �����������������������������U����   SVW��@����0   �������E�Q����B(�H�у�;�衯���E�     _^[���   ;�舯����]��������������������������������������U����   SVW��@����0   �������E�Q����B(�H�у�;��!����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B,�H�у�;�衮���E�     _^[���   ;�舮����]��������������������������������������U����   SVW��@����0   �������E�Q����B,�H0�у�;��!����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;�蠭���E�     _^[���   ;�臭����]�������������������������������������U����   SVW��@����0   �������EP����Q$�B\�Ѓ�;��#���_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP����Q�B �Ѓ�;�賬��_^[���   ;�裬����]���������������������������������U����   SVW��@����0   �������EP�MQ����B�H(�у�;��?���_^[���   ;��/�����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B��  �у�;������_^[���   ;�谫����]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H�Q�҃�;��L���_^[���   ;��<�����]��������������������������U����   SVW��@����0   �������EP����Q�B�Ѓ�;�����_^[���   ;��Ӫ����]���������������������������������U���  SVW�������E   ������E�P�M�]����M��l����uǅ����    �M���q���������   j�E�P芞������u*�E�P�|�������uǅ����    �M��q���������Tj�EP�N�������u*�EP��������uǅ���    �M��Hq��������ǅ���   �M��.q�������R��P�x�
�h���XZ_^[��  ;�諩����]�   ��
����   ��
parent �����������������������������������������������������������������������������U����   SVW��@����0   �������EP�MQ����B�H�у�;������_^[���   ;�������]�����������������������������U����   SVW��@����0   �������EP����Q��  �Ѓ�;�萨��_^[���   ;�耨����]������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��   �Ѓ�;�����_^[���   ;�������]����������������������������������U����   SVW��@����0   �������EP�MQ����B�H�у�;�蟧��_^[���   ;�菧����]�����������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��,���_^[���   ;�������]��������������������������U����   SVW��@����0   �������EP�MQ����B�H�у�;�迦��_^[���   ;�详����]�����������������������������U����   SVW��@����0   �������EP�MQ�UR����H��  �҃�;��I���_^[���   ;��9�����]�����������������������U����   SVW������9   �������EP�� ���Q����B���  �у�;��٥��P�M�X����� ����!m���E_^[���   ;�貥����]��������������������������������U����   SVW��@����0   �������EP����Q��L  �Ѓ�;��P���_^[���   ;��@�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H��D  �҃�;��٤��_^[���   ;��ɤ����]�����������������������U���$  SVW�������I   ������ǅ8���    �=�� t!������P����D�����8����������������O����8���������������������������R�M貭����8�����t��8����������ik����8�����t��8�����������Lk���E_^[��$  ;��ݣ����]�����������������������������������������������������������U����   SVW������9   ������� ���P����Q���  �Ѓ�;��]���P�M�ܬ���� ����j���E_^[���   ;��6�����]������������������������������������U����   SVW������9   ������� ���P����Q�B$�Ѓ�;��Т��P�M�O����� ����j���E_^[���   ;�詢����]���������������������������������������U����   SVW��@����0   ������j�EP�y������E_^[���   ;��@�����]������������������������������U����   SVW��@����0   �������EP�MQ�UR����H�Q�҃�;��ܡ��_^[���   ;��̡����]��������������������������U����   SVW��@����0   �������EP�MQ�UR����H��H  �҃�;��i���_^[���   ;��Y�����]�����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bd��;������_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q$�B`�Ѓ�;�肠��_^[���   ;��r�����]� �����������������������������U����   SVWQ������<   ������Y�M���E�P�����Q����B$�H �у�;�����P�M膩��������Og���E_^[���   ;��������]� �������������������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��p���_^[���   ;��`�����]������������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B0��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;�萞��_^[���   ;�耞����]������������������������������U����   SVWQ������<   ������Y�M���E�P�����Q����B$�H$�у�;�����P�M薧��������_e���E_^[���   ;�������]� �������������������������������������������U����   SVWQ������<   ������Y�M��EP�����Q�M��W�����耮���������d���E_^[���   ;��d�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B,�M��P��;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;�耜��_^[���   ;��p�����]������������������������������U����   SVWQ������<   ������Y�M������P����Q,�M��B��;�����P�M芥��������Sc���E_^[���   ;�������]� �������������������������������U����   SVWQ������<   ������Y�M������P����Q,�M��B<��;��{���P�M������������b���E_^[���   ;��T�����]� �������������������������������U����   SVWQ��4����3   ������Y�M�����P$��M��Bp��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B,��;�胚��_^[���   ;��s�����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B8��;�裙��_^[���   ;�蓙����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P(��M��B(��;��3���_^[���   ;��#�����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B��;��Ø��_^[���   ;�賘����]���������������������������������U����   SVWQ������9   ������Y�M���E�P�� ���Q����B$�H�у�;��G���P�M��t���� ����K����E_^[���   ;�� �����]� �������������������������������������������U����   SVWQ������9   ������Y�M���EP�� ���Q����B,�M��P@��;�觗��P�M�+t���� �������E_^[���   ;�耗����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H,�Q�҃�;�����_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B4��;�蓖��_^[���   ;�胖����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B(��;��#���_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B��;�賕��_^[���   ;�裕����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B ��;��C���_^[���   ;��3�����]���������������������������������U����   SVWQ��4����3   ������Y�M�����P,��M��B$��;��Ӕ��_^[���   ;��Ô����]���������������������������������U����   SVWQ��4����3   ������Y�M���E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP����Q(�M����   ��;��7���_^[���   ;��'�����]�( ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR����P(�M��B��;�諓��_^[���   ;�蛓����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����;��#���_^[���   ;�������]� ������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����   ��;�蟒��_^[���   ;�菒����]� ��������������������������U����   SVWQ��$����7   ������Y�M��E�P�M��Z����u3��.�E��tǅ$���   �
ǅ$���    �M��$�����   R��P�<�
覥��XZ_^[���   ;�������]�    D�
����   P�
c ����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��[���_^[���   ;��K�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P(�M��B��;�����_^[���   ;��א����]� ����������������������������������U����   SVWQ��0����4   ������Y�M��} t2��EP�M�Q����B �H$�у�;��d�����tǅ0���   �
ǅ0���    ��0���_^[���   ;��4�����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�UR����H �QL�҃�;�跏��_^[���   ;�觏����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��BX��;��>���_^[���   ;��.�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B`��;��Ύ��_^[���   ;�辎����]� �������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��`���_^[���   ;��P�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;�����_^[���   ;��׍����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;��g���_^[���   ;��W�����]� ����������������������������������U����   SVWQ������?   ������Y�M��M��ǒ���E�P�M��[����uǅ���    �M���t��������$�E�P�M�P��ǅ���   �M���t�������R��P���
�R���XZ_^[���   ;�蕌����]�    ��
����   ��
str ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;������_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��  �у�;�臋��_^[���   ;��w�����]� ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B���   �у�;�� ���_^[���   ;��������]������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�苊��_^[���   ;��{�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bx��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�諉��_^[���   ;�蛉����]� ����������������������U����   SVWQ��0����4   ������Y�M��EP�M��ӗ����tE�M��Q�M��������t2�U��0R�M�譗����t�E��HP�M�蚗����tǅ0���   �
ǅ0���    ��0���_^[���   ;�������]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��k���_^[���   ;��[�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bt��;������_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�苇��_^[���   ;��{�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M���  ��;�諆��_^[���   ;�蛆����]� ����������������������U����   SVWQ��0����4   ������Y�M��EP�M�蜅����t2�M��Q�M�艅����t�U��R�M��v�����tǅ0���   �
ǅ0���    ��0���_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�苅��_^[���   ;��{�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bh��;�����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bp��;�讄��_^[���   ;�螄����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��;���_^[���   ;��+�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;��ǃ��_^[���   ;�跃����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bx��;��N���_^[���   ;��>�����]� �������������������������U����   SVWQ��0����4   ������Y�M��EP�M��S����tE�M��Q�M���R����t2�U��R�M���R����t�E��$P�M���R����tǅ0���   �
ǅ0���    ��0���_^[���   ;�臂����]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�����_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bp��;�螁��_^[���   ;�莁����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B|��;��.���_^[���   ;�������]� �������������������������U����   SVWQ��0����4   ������Y�M��EP�M��aJ����t2�M��Q�M��NJ����t�U��R�M��;J����tǅ0���   �
ǅ0���    ��0���_^[���   ;��z�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;�����_^[���   ;�������]� ����������������������U����   SVWQ������?   ������Y�M��E�    �E�    �E�P�M��)�����u3���   �}� u)������I���P�M�k��������g���   �   ��h0`����P�M�Q����B���   �у�;��9���E��}� uj��M��/���3��Lj �E�P�M�Q�M��
g����u�E�P�|L����3��&j �E��P�M�Q�M�����E�P�WL�����   R��P�p�
�r���XZ_^[���   ;��~����]�    x�
����   ��
����   ��
c len ������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;���}��_^[���   ;���}����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��{}��_^[���   ;��k}����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B\��;��}��_^[���   ;���|����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bd��;��|��_^[���   ;��|����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bl��;��.|��_^[���   ;��|����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bt��;��{��_^[���   ;��{����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��Bd��;��N{��_^[���   ;��>{����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bl��;���z��_^[���   ;���z����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��kz��_^[���   ;��[z����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;���y��_^[���   ;���y����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B`��;��y��_^[���   ;��~y����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bh��;��y��_^[���   ;��y����]� �������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��x��_^[���   ;��x����]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P(�M��B$��;��7x��_^[���   ;��'x����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q�B�Ѓ�;��w��_^[���   ;��w����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H4�у�;��:w��_^[���   ;��*w����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B4��;��v��_^[���   ;��v����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��Kv��_^[���   ;��;v����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H8�у�;���u��_^[���   ;���u����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q$�M��Bl��;��^u��_^[���   ;��Nu����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H$�QP�҃�;���t��_^[���   ;���t����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�HT�у�;��jt��_^[���   ;��Zt����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��B��;���s��_^[���   ;���s����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H�у�;��zs��_^[���   ;��js����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B$�H,�у�;���r��_^[���   ;���r����]� �������������������������������������U����   SVW��@����0   �������EP�MQ����B���  �у�;��|r��_^[���   ;��lr����]��������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��r��_^[���   ;�� r����]������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��q��_^[���   ;��q����]� ����������������������U����   SVWQ��4����3   ������Y�M���j�EP�MQ����B(�M��P��;��(q��_^[���   ;��q����]� �����������������������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��p��_^[���   ;��p����]�����������������������U����   SVW��@����0   �������EP�MQ�UR����H���  �҃�;��9p��_^[���   ;��)p����]�����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����   ��;��o��_^[���   ;��o����]� ��������������������������U����   SVWQ��0����4   ������Y�M��} t	ƅ3����ƅ3��� ��3���P�M���y��_^[���   ;��6o����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B,��;���n��_^[���   ;��n����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B(�M��P ��;��Zn��_^[���   ;��Jn����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��} u3��'��EP�M�Q����B �H(�у�;���m���   _^[���   ;��m����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��B8��;��Mm��_^[���   ;��=m����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;���l��_^[���   ;���l����]� ������������������������U����   SVWQ��4����3   ������Y�M�����P��M����   ��;��pl��_^[���   ;��`l����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;���k��_^[���   ;���k����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BT��;��~k��_^[���   ;��nk����]� �������������������������U����   SVWQ������<   ������Y�M��� ���P�M�|��P�M��&J��������� ����S�������_^[���   ;���j����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BP��;��~j��_^[���   ;��nj����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��  �у�;��j��_^[���   ;���i����]� ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q��   �Ѓ�;��i��_^[���   ;��ti����]����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M����   ��;���h��_^[���   ;���h����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B(�M��P|��;��h��_^[���   ;��zh����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��P\��;��
h��_^[���   ;���g����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��s����tE�M��Q�M���r����t2�U��0R�M���r����t�E��HP�M���r����tǅ0���   �
ǅ0���    ��0���_^[���   ;��7g����]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BH��;��f��_^[���   ;��f����]� �������������������������U����   SVWQ��4����3   ������Y�M�����E�$����P(�M��BT��;��Ff��_^[���   ;��6f����]� ���������������������������������U����   SVWQ��4����3   ������Y�M�����E�$����P�M��B(��;���e��_^[���   ;��e����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M���  ��;��Ge��_^[���   ;��7e����]� ����������������������������������U����   SVWQ��0����4   ������Y�M��E��� �$�M��y����tD�M���A�$�M��y����t(�U���B�$�M��~y����tǅ0���   �
ǅ0���    ��0���_^[���   ;��md����]� ��������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B<��;���c��_^[���   ;���c����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��BH��;��~c��_^[���   ;��nc����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B��;��c��_^[���   ;���b����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B@��;��b��_^[���   ;��b����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��PX��;��*b��_^[���   ;��b����]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$����P�M��B ��;��a��_^[���   ;��a����]� ���������������������������������U����   SVWQ��0����4   ������Y�M��EP�M��/����tE�M��Q�M��}/����t2�U��R�M��j/����t�E��$P�M��W/����tǅ0���   �
ǅ0���    ��0���_^[���   ;���`����]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BD��;��^`��_^[���   ;��N`����]� �������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$����P(�M��BP��;���_��_^[���   ;���_����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���Q�E�$����P�M��B$��;��h_��_^[���   ;��X_����]� �����������������������������������U����   SVWQ��0����4   ������Y�M��EQ� �$�M���<����t@�MQ�A�$�M���<����t&�UQ�B�$�M��<����tǅ0���   �
ǅ0���    ��0���_^[���   ;��^����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B8��;��^��_^[���   ;��^����]� �������������������������U����   SVWQ������=   ������Y�M�j �M�U�����E���h0`����P�M�Q����B���   �у�;��]���Eԃ}� uj��M��^��3��dj �E�P�M�Q�M�_b���E�P�M��G����t �M�Q�U�R�M��d����tǅ���   �
ǅ���    ������E�E�P�*�����E�R��P�4�p��XZ_^[���   ;���\����]�    <����   Hmem ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��BL��;��>\��_^[���   ;��.\����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B0��;���[��_^[���   ;��[����]� �������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��B<��;��][��_^[���   ;��M[����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;���Z��_^[���   ;���Z����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP����Q(�M��BL��;��~Z��_^[���   ;��nZ����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B��;��Z��_^[���   ;���Y����]� �������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��BD��;��Y��_^[���   ;��Y����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;��-Y��_^[���   ;��Y����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��B4��;��X��_^[���   ;��X����]� �������������������������U����   SVWQ��4����3   ������Y�M����EP����Q(�M��B@��;��MX��_^[���   ;��=X����]� ������������������������U����   SVWQ��4����3   ������Y�M����EP����Q�M��B��;���W��_^[���   ;���W����]� ������������������������U����   SVWQ��4����3   ������Y�M���EPj�����Q�M��B��;��lW���E�_^[���   ;��YW����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���j �EP����Q�M��B��;���V���E�_^[���   ;���V����]� ������������������������������������U����   SVWQ��4����3   ������Y�M���j j�����P�M��B��;��oV���E�_^[���   ;��\V����]��������������������������U����   SVWQ��4����3   ������Y�M��M��4c��_^[���   ;��V����]������������������U����   SVWQ��4����3   ������Y�M�j j �E�P�M�i!���E�_^[���   ;��U����]� ��������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�H�у�;��JU��_^[���   ;��:U����]� �������������������������������������U����   SVWQ��0����4   ������Y�M���EP�M�Q����B�H�у�;���T����uǅ0���   �
ǅ0���    ��0���_^[���   ;��T����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M����   ��;��$T��_^[���   ;��T����]� �������������������������������U����   SVWQ��4����3   ������Y�M�����P��M��B��;��S��_^[���   ;��S����]���������������������������������U����   SVWQ��(����6   ������Y�M��EP�M��-:���E�M��:E��_^[���   ;��5S����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BX�Ѓ�;���R��_^[���   ;��R����]�������������������������U����   SVWQ��(����6   ������Y�M��EP�M��M9���E�EP�M���9��_^[���   ;��QR����]� ����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q������   �H`�у�;���Q��_^[���   ;���Q����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M��Bt��;��nQ��_^[���   ;��^Q����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P�M��Bl��;���P��_^[���   ;���P����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�hF  �EP�MQ�M���a��_^[���   ;��wP����]� ����������������������������������U����   SVWQ��4����3   ������Y�M�h#  �EP�MQ�M��Va��_^[���   ;��P����]� ����������������������������������U����   SVWQ��(����6   ������Y�M���EP����Q�M����   ��;��O���E�}� u3���M��&��_^[���   ;��vO����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �B�Ѓ�;��O��_^[���   ;���N����]�������������������������U����   SVWQ��4����3   ������Y�M���EP����Q�M����   ��;��N��_^[���   ;��N����]� ����������������������U���  SVWQ��X����j   ������Y�M��-���M���E��8 u��   �EP��l����8��j h|`�������B*��P�������8��j j���l���Q������R������P�9����P������Q�G����P�����R�G����P�E��������tǅX���   �
ǅX���    ��X�����c�������������������������������������������������v5����l��������c�����t�E�P�N�����E�_^[�Ĩ  ;��)M����]� ������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�D�����M���E�_^[���   ;��L����]� �������������������U����   SVWQ��4����3   ������Y�M��E�P�R����_^[���   ;��0L����]����������������̋�`��`��`��`��`��`��` ��`$��`(��`,��`0��`4��`8��`<��`@��`�������������U����   SVW��@����0   ������EP�M���   Q�UR�8����_^[���   ;��wK����]���������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVW��@����0   ������E�M�H4�E�@d�E�@8�J�E�@<�J�E�@@�D�E�@D+^�E�@H�\�E�@L#\�E�@P�s�E�@l1]�E�@X�\�E�@\�]�E�@`&^�E�@d]�E�@T]�E�@h�t�E�@p�]�E�@t	]�E�M�H �E�M��E�M�H0�E�M�H(�E�@,    _^[��]����������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�_^[��]� ��������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U���h  SVW�������Z   ������j h�   ��\���P������j �EP�MQ�UR�EP��\���Q�"�����E �E�h�   ��\���P�MQ�URj�����R��P����Y��XZ_^[��h  ;��5F����]Ë�   �\����   np ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M���1���M���E�_^[���   ;���D����]�����������������������������U����   SVWQ��4����3   ������Y�M��E��x^� �E���`�@�E�_^[��]���������������������U����   SVWQ��4����3   ������Y�M��E��M��E��@    �E��@    �E�_^[��]� ���������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q������   �H,�у�;��C���E�_^[���   ;��C����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    ��EP�M�Q������   �H(�у�;��C���E�_^[���   ;���B����]� ��������������������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��M�H�E�_^[��]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��    �E��E�@�E�_^[��]� ���������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E�P�uD�����E��     _^[���   ;��A����]���������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVW��@����0   ������EE_^[��]����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL��  �у�;��'@��_^[���   ;��@����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL�QT�҃�;��?��_^[���   ;��?����]� ����������������������������������U����   SVW��@����0   �����󫡸����   �􋑈   ��;��5?��_^[���   ;��%?����]�����������������������������������U����   SVW��@����0   �����󫡸��HL��Q��;���>��_^[���   ;��>����]�������������������������U����   SVW��@����0   �����󫡸��HL���   ��;��h>��_^[���   ;��X>����]����������������������U����   SVW��@����0   �����󫡸��HL����;��>��_^[���   ;���=����]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL�B\�Ѓ�;��=��_^[���   ;��=����]� �����������������������������U����   SVW��@����0   �����󫡸��HL��  ��;��(=��_^[���   ;��=����]����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL��   �Ѓ�;��<��_^[���   ;��<����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M��B��;��4<��_^[���   ;��$<����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�BX�Ѓ�;��;��_^[���   ;��;����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL���   �у�;��G;��_^[���   ;��7;����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�BP�Ѓ�;���:��_^[���   ;��:����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ����BL�M���H  ��;��K:��_^[���   ;��;:����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;���9��_^[���   ;��9����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;��[9��_^[���   ;��K9����]�������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;���8���E�     _^[���   ;���8����]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��q8���E�     _^[���   ;��X8����]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;���7���E�     _^[���   ;���7����]��������������������������������������U���0  SVWQ�������L   ������Y�M��M������h�  �������)��P��������*��j �E�P������Q�M��Y�����uǅ����   �
ǅ����    �������������������4����������tǅ���    �M������������M����������M���������R��P�d)�}J��XZ_^[��0  ;���6����]Ð   l)����   x)dat ��������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B`�Ѓ�;��6��_^[���   ;��6����]����������������������������U����   SVW��@����0   �����󫡸��H�􋑘   ��;��5��_^[���   ;��5����]����������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B4�Ѓ�;��N5��_^[���   ;��>5����]����������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M����   ��;���4��_^[���   ;���4����]� ����������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B0�Ѓ�;��n4��_^[���   ;��^4����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;���3��_^[���   ;���3����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����QL�M���l  ��;��o3��_^[���   ;��_3����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;���2��_^[���   ;���2����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B,�Ѓ�;��~2��_^[���   ;��n2����]����������������������������U����   SVWQ��4����3   ������Y�M���j �E�P����QL�B8�Ѓ�;��2��_^[���   ;���1����]��������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M����   ��;��1��_^[���   ;��1����]� ����������������������U����   SVWQ������:   ������Y�M���EP�M�Q�����R����HL��  �҃�;��!1��P�M�/��������]����E_^[���   ;���0����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL�Hh�у�;��0��_^[���   ;��z0����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL��D  �Ѓ�;��0��_^[���   ;���/����]�������������������������U���0  SVWQ�������L   ������Y�M��M������h�  �������5!��P�������#��j �E�P������Q�M�������uǅ����   �
ǅ����    ��������������������,����������tǅ���    �M�����������M�����������M����������R��P�41�B��XZ_^[��0  ;���.����]Ð   <1����   H1dat ��������������������������������������������������������������������U����   SVWQ������:   ������Y�M���EP�M�Q�����R����HL�Q�҃�;��D.��P�M�8,������������E_^[���   ;��.����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M���p  ��;��-��_^[���   ;��-����]� ����������������������������������U���  SVWQ�������F   ������Y�M��M�����h�  ���������P������� ��j �E�P������Q�M�������uǅ����   �
ǅ����    �������������������l*����������t�M�����M��	���E��M�����P�M�96���M��|	���ER��P��3�B@��XZ_^[��  ;��,����]�    �3����   �3dat ������������������������������������������������������������������������U���  SVWQ�������F   ������Y�M��M��<���h�  ������u��P�������D��j �E�P������Q�M��������uǅ����   �
ǅ����    �������������������)����������t�M�|���M��J���E��M����P�M��4���M��,���ER��P��4��>��XZ_^[��  ;��5+����]�    �4����   5dat ������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BL�Ѓ�;��*��_^[���   ;��{*����]�������������������������U����   SVW��@����0   �����󫡸��H�􋑜   ��;��(*��_^[���   ;��*����]����������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;��)��_^[���   ;��)����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL��(  �Ѓ�;��K)��_^[���   ;��;)����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;���(��_^[���   ;���(����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�B�Ѓ�;��n(��_^[���   ;��^(����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;���'��_^[���   ;���'����]�������������������������U���0  SVWQ�������L   ������Y�M��M������h�  �������%��P����������j �E�P������Q�M��y�����uǅ����   �
ǅ����    ��������������������$����������tǅ���    �M������������M�����������M����������R��P�D9�:��XZ_^[��0  ;���&����]Ð   L9����   X9dat ��������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;��;&��_^[���   ;��+&����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL�Q@�҃�;���%��_^[���   ;��%����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M����  ��;��K%��_^[���   ;��;%����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP������   �M����   ��;���$��_^[���   ;���$����]� �����������������������������������U���8  SVWQ�������N   ������Y�M��M�����h�  ����������P����������j �E�P������Q�M��I�����uǅ����   �
ǅ����    �������������������!����������t �x^�� ����M��� ��݅ �����M��L ��ݝ����M�� ��݅���R��P�|<�g7��XZ_^[��8  ;��#����]ÍI    �<����   �<dat ����������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL���   �Ѓ�;���"��_^[���   ;���"����]�������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��BP��;��"��_^[���   ;��"����]������������������������������U���  SVWQ�������F   ������Y�M��M��|���h�  ��������P���������j �E�P������Q�M��	�����uǅ����   �
ǅ����    �������������������\����������t�M��&���M������E�,�M��#����M���P�Q�P�Q�@�A�M��\����ER��P��>�"5��XZ_^[��  ;��e!����]�    �>����   �>dat ������������������������������������������������������������������������U���  SVWQ�������F   ������Y�M��M�����h�  ������U��P�������$��j �E�P������Q�M�������uǅ����   �
ǅ����    ������������������������������t�M�n%���M��*����E�,�M�������M���P�Q�P�Q�@�A�M�������ER��P� @��3��XZ_^[��  ;�� ����]�    (@����   4@dat ������������������������������������������������������������������������U���  SVWQ�������F   ������Y�M��M�����h�  ���������P����������j �E�P������Q�M��I�����uǅ����   �
ǅ����    �����������������������������t�M�$���M�������E�,�M��c����M���P�Q�P�Q�@�A�M������ER��P��A�b2��XZ_^[��  ;������]�    �A����   �Adat ������������������������������������������������������������������������U���  SVWQ�������F   ������Y�M��M��\���h�  ��������P�������d��j �E�P������Q�M��������uǅ����   �
ǅ����    �������������������<����������t�M�"���M��j����E�,�M������M���P�Q�P�Q�@�A�M��<����ER��P��B�1��XZ_^[��  ;��E����]�    �B����   �Bdat ������������������������������������������������������������������������U���0  SVWQ�������L   ������Y�M��M������h�  �������5��P���������j �E�P������Q�M�������uǅ����   �
ǅ����    ������������������������������tǅ���    �M������������M������������M�����������R��P�4D�/��XZ_^[��0  ;�������]Ð   <D����   HDdat ��������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��B(��;��P��_^[���   ;��@����]������������������������������U����   SVWQ��4����3   ������Y�M�����PL��M���L  ��;�����_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �B<�Ѓ�;��k��_^[���   ;��[����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL��  �҃�;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�Bd�Ѓ�;��~��_^[���   ;��n����]����������������������������U���0  SVWQ�������L   ������Y�M��M��l���h�  �������
��P�������t��j �E�P������Q�M��������uǅ����   �
ǅ����    �������������������L����������tǅ���    �M��x����������M��Z���������M��Z��������R��P��G�,��XZ_^[��0  ;��`����]Ð   �G����   �Gdat ��������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M����   ��;����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL���   �у�;��G��_^[���   ;��7����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�Bl�Ѓ�;�����_^[���   ;������]����������������������������U���  SVWQ�������F   ������Y�M��M�����h�  ���������P��������	��j �E�P������Q�M��I�����uǅ����   �
ǅ����    �����������������������������t�M����M�������E�,�M��c����M���P�Q�P�Q�@�A�M������ER��P��J�b)��XZ_^[��  ;������]�    �J����   �Jdat ������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P������   �BP�Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ������9   ������Y�M���j �EP�M�Q�� ���R����HL���   �҃�;�����M���P�Q�P�Q�@�A�E_^[���   ;��S����]� ����������������������������������������������U����   SVWQ������9   ������Y�M���j�EP�M�Q�� ���R����HL���   �҃�;������M���P�Q�P�Q�@�A�E_^[���   ;������]� ����������������������������������������������U����   SVW��@����0   ������E���M���;��<��_^[���   ;��,����]��������������������������U����   SVW��@����0   �������EP�MQ�U��M�P��;�����_^[���   ;�������]���������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�M��M�B��;��[��_^[���   ;��K����]�������������������������U����   SVW��@����0   �������EP�M��M�B��;�����_^[���   ;�������]���������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����HL���   �҃�;��x��_^[���   ;��h����]� �����������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;�� ��_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��B<��;����_^[���   ;��{����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL�B$�Ѓ�;����_^[���   ;������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL��,  �҃�;����_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����BL�H(�у�;����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL�B �Ѓ�;����_^[���   ;������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL��4  �у�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��BH��;����_^[���   ;������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL���   �҃�;��$��_^[���   ;������]� �������������������������������U����   SVWQ��(����6   ������Y�M���E�P����QL���   �Ѓ�;�����E�}� u)��j �EP�M�Q����BL���   �у�;��{����M��!��P�M�����_^[���   ;��X����]� ���������������������������������������������������U���  SVW�������B   ������M��d����M��}���} t�M��Y�����u"ǅ����   �M�������M�������������Qj�M��)���P�M� ���M������E�E�E��E�Ph<��������������M��t����M����������R��P��T���XZ_^[��  ;��K����]�   �T����   �T����   �Tactive mu ������������������������������������������������������������������������������U���  SVW�������B   ������M������M��-���} t�M��	�����u"ǅ����   �M��w����M������������Qj�M������P�M�c���M�������E�E�E��E�Ph=���M�����������M��$����M��I��������R��P�(V���XZ_^[��  ;���	����]�   0V����   OV����   HVactive mu ������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�����PL��M����  ��;��@	��_^[���   ;��0	����]������������������������������U����   SVWQ��$����7   ������Y�M��M�������E�}�t�}�t�}�tǅ$���    �
ǅ$���   ��$���_^[���   ;������]���������������������������������U����   SVW��@����0   �������EP�MQ����BL���   �у�;��<��_^[���   ;��,����]��������������������������U����   SVW��@����0   �������E�Q����B���   �у�;������E�     _^[���   ;������]�����������������������������������U����   SVW��4����3   �������+���E��}� u3��a��j �EP�MQ�UR�E�P����Q��h  �Ѓ�;��0����u+�}� t��E�P����Q@�B�Ѓ�;�����E�    �E�_^[���   ;�������]��������������������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;����_^[���   ;��p����]������������������������������U����   SVW��@����0   �������j �EPj �MQ������P�UR�EP����Q��h  �Ѓ�;�����_^[���   ;�������]�������������������������������������U���T  SVWQ�������U   ������Y�M��V ���E�}� u3��  �E�    �E�    �E�    �M������M�������E�E��E��E��EPh]  �M������j j �E�P�M��������u��   �M�����E���E��Eȃ}� ��   �M������E��EȉE��E�Ph�   ��������u�   �}� u�~j �M��N����Eԃ}� u�i�E�P�M��&����E�P������}� t��E�P����Q@�B�Ѓ�;�����E�    �`����E쉅�����M������M������������W�}� t��E�P����Q@�B�Ѓ�;��:���E�    �E�P�|����ǅ����    �M��<����M��]���������R��P�@\���XZ_^[��T  ;�������]� �   H\����   c\����   `\cd ctr �����������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QL���   �Ѓ�;�����_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����BL��   �у�;��[��_^[���   ;��K����]� ��������������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����Q���   �Ѓ�;�����_^[���   ;������]��������������������������������������U����   SVWQ��4����3   ������Y�M��E��M�H�E��M$�H��h�MhMh�Mh�L�E��HQ�U R�EP�MQ���E�$�UR�E��HQ�U�R����HL���   �҃�4;��� ��_^[���   ;��� ����]�  ������������������������������������������������������U����   SVW��@����0   �������EP�MQ�UR����HL���   �҃�;��i ��_^[���   ;��Y ����]�����������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q���   �Ѓ�;������_^[���   ;��������]����������������������������������U����   SVWQ��4����3   ������Y�M���j �EP�M�Q����BL�HD�у�;��x���_^[���   ;��h�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�M�Q����BL�HD�у�;������_^[���   ;��������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j �EP�M�Q����BL�HH�у�;��x���_^[���   ;��h�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���j�EP�M�Q����BL�HH�у�;������_^[���   ;��������]� �����������������������������������U���  SVWQ�������B   ������Y�M��EP����������h�  ��$�������P����������j������Q�����R�M��3�����������������������_^[��  ;��3�����]� ����������������������������������������������U����   SVW��@����0   �������EP����Q���   �Ѓ�;������_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;��G���_^[���   ;��7�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;������_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL�H<�у�;��J���_^[���   ;��:�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;������_^[���   ;�������]� ����������������������������������U���  SVWQ�������B   ������Y�M�j����������h�  ��$��������P���������j������P�����Q�M�������������������������_^[��  ;�������]���������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HL�Q�҃�;�����_^[���   ;��w�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M���t  ��;�����_^[���   ;��������]� ����������������������������������U���  SVWQ�������B   ������Y�M��EP�����������h�  ��$�������P����������j������Q�����R�M��C��������������������&���_^[��  ;��C�����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP����������h�  ��$����^���P������-���j������Q�����R�M�胾��������(����������f���_^[��  ;�������]� ����������������������������������������������U����   SVW��@����0   �������EP�MQ����BL���   �у�;�����_^[���   ;��������]��������������������������U���  SVWQ�������B   ������Y�M��EP�������&���h�  ��$����.���P����������j������Q�����R�M��S��������������������6���_^[��  ;��S�����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����  ��;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����  ��;��W���_^[���   ;��G�����]� ����������������������������������U���  SVWQ�������B   ������Y�M����E�$����������h�  ��$����e���P������4���j������P�����Q�M�芻��������/����������m���_^[��  ;�������]� �����������������������������������������������������U���  SVWQ�������B   ������Y�M��EP�������M���h�  ��$�������P������m���j������Q�����R�M��ú��������h�������������_^[��  ;��������]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP����������h�  ��$��������P���������j������Q�����R�M�������������������������_^[��  ;�������]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP�����������h�  ��$�������P����������j������Q�����R�M��C��������������������&���_^[��  ;��C�����]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP����������h�  ��$����^���P������-���j������Q�����R�M�胸��������(����������f���_^[��  ;�������]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP����������h�  ��$�������P������m���j������Q�����R�M��÷��������h�������������_^[��  ;��������]� ����������������������������������������������U���  SVWQ�������B   ������Y�M��EP����������h�  ��$��������P���������j������Q�����R�M�������������������������_^[��  ;�������]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BL���   �у�;�����_^[���   ;��w�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����BL�M����   ��;�����_^[���   ;��������]� ����������������������������������U���  SVWQ�������B   ������Y�M��EP�����������h�  ��$�������P����������j������Q�����R�M��C��������������������&���_^[��  ;��C�����]� ����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M���P  ��;������_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���E�P����QL�BL�Ѓ�;��^���_^[���   ;��N�����]����������������������������U����   SVW��@����0   �����󫡸��HL��@  ��;������_^[���   ;��������]����������������������U����   SVWQ��4����3   ������Y�M���EP����QL�M���T  ��;�����_^[���   ;��{�����]� ����������������������U����   SVW��@����0   ������E;Et�&�} t �} t�} t�EP�MQ�UR�Ⱥ����_^[���   ;�������]�������������������������������U����   SVW��@����0   ������E;Et�&�} t �} t�} t�EP�MQ�UR�H�����_^[���   ;�������]�������������������������������U����   SVWQ��4����3   ������Y�M��M�������E�� �`�E�_^[���   ;�������]����������������������U����   SVWQ��4����3   ������Y�M��E�� �`�E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E�� �`�E��@    �E�_^[��]�����������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��4����3   ������Y�M��E��     �E�_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��E�� �`��E��HQ����Bl�H�у�;�����_^[���   ;��r�����]��������������������������������U����   SVWQ��4����3   ������Y�M�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M���j�E��Q����BH��|  �у�;������_^[���   ;�������]�������������������������������������U����   SVWQ��4����3   ������Y�M��M��3����E��t�E�P�!������E�_^[���   ;��=�����]� ������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ�UR����HH���   �҃�;������_^[���   ;��������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���   �҃�;��T���_^[���   ;��D�����]� �������������������������������U����   SVW��@����0   �������EP����QH��Ѓ�;������_^[���   ;��������]����������������������������������U����   SVW��@����0   �������h�  ����HH��҃�;��t���_^[���   ;��d�����]����������������������������������U����   SVW��4����3   ������h  ��������E��}� u3��tj �EPh�  �M��������u�.�,j �EPh(  �M��������u��j j�M������E��-�}� t��E�P����Q@�B�Ѓ�;������E�    3�_^[���   ;�������]�������������������������������������������������U����   SVW��@����0   �����󫡸��HH���  ��;�����_^[���   ;�������]����������������������U����   SVW��4����3   ������h�  �������E��}� u3��B�EP�MQ�M�������u+�}� t��E�P����Q@�B�Ѓ�;������E�    �E�_^[���   ;��e�����]���������������������������������������������������U����   SVW��@����0   �����󫡸��HH��  ��;������_^[���   ;��������]����������������������U����   SVW��@����0   �������EP�MQ����BH�H�у�;�����_^[���   ;�������]�����������������������������U����   SVW��@����0   �������*E�YE�X0a�,��E�EP�MQ�UR������_^[���   ;�������]����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;�����_^[���   ;�������]� ����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����BH��0  �у�;�����_^[���   ;�� �����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;�����_^[���   ;�������]� ����������������������������������U����   SVW��@����0   �������EP�MQ����BH���  �у�;�����_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M��E�M� +_^[��]� ��������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;��[���_^[���   ;��K�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����HH���  �҃�;������_^[���   ;��������]� �����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;��[���_^[���   ;��K�����]�������������������������U����   SVW��@����0   ��������E�$���E�$���x^�$�EP�M�W������$腬�����$�MQ�M�����_^[���   ;�������]��������������������������������������������U���   SVW�������H   �����󫍍���������P�EP�M�Q�M�������E�$���E�$���E��$�Ϋ�����$���E�$���E�$���E��$蜫�����$���E�$���E�$���E��$�j������$����������P�EP�M����R��P����3���XZ_^[��   ;��v�����]ÍI    ������   Ăv ��������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���j �E��Q����BH��|  �у�;������_^[���   ;�������]�������������������������������������U���D  SVW��������   ������M�����E��E�    �M�f����E��E�    �E�    �E�    �E�    �}� u
�   ��  �M�~���=�  �  j h:  �M������E��M������E�ǅP���    �M������,����M莞���� ����M�������������������E�    �	�E����E��E�;E���   �� ��� ��   j��E�P�� ����g�����t�����t����tek�t��������N���9E�t�k�t��������w���������������;�P���~��������P���k�t�����������EԉE��6�E����M�����,�����,����D;Du�Eԃ��E��	�Eԃ��E������}� tj �EP�M�������u
�%  �   �}� tz�M��������tn�M��C���;E�ua��h�`� ���%PkM�Q����B���  �у�;��]����E��}� u
��  �  �E�PkM�Q�U�R�M�����P��������h�`� ���)PkM�Q����B���  �у�;�������E��}� u
�b  �]  �E�PkM�Q�U�R�E�P�=�������P��� ~K��h�`� ���.P��P�������Q����B���   �у�;������E��}� u
��  ��  j��E�P�M跩����u
��  ��  �}� tj�EP�M�裠����u
�  �  �}� t�M������������
ǅ����    �������E��M�����E��E�    �E�    �	�E����E��E�;E���  �� ��� ��  j��E�P�� ���豲����t�����t������  k�t�������蔯��9E�t�k�t��������_���������ǅ����    ǅ\���    ǅh���    ���h�������h���k�t�����������9�h�����  ��h���Pk�t��������u�����u봋�h���Pk�t��������������D�����D�������\����U���,��������\�������\�����D�������\����U�����\�������\�����D�������\����U���,����D����\�������\�����D�����   ��\����E�����\�������\�����D�������\����U���,����D����\�������\�����D�����   ��\����E�����\�������\�����D�������\����U���,����D����\�������\�����D�����   ��\����E�����\�������\����=�����\��������������� �v  j�������+���P�E�P�����詗��ǅ\���    ������;�����|6ha� ���ZPh�`hL[�C�����h�`� ���ZP������������;�����|
�}	  �x	  ��\����M����������}� t3k�����E�kM�M����P�Q�P�Q�P�Q�P�Q�@�Ak�����E�kM�Mȋ��P�Q�P�Q�P�Q�P�Q�@�A��\���;�������   ��\����M���;�������   ��\����M��D���������D�����\����M��T�����8�����8���������������wj�������$�P���D�������,����Uԉ�F��D�������,����UԉT�.��D�������,����UԉT���D�������,����UԉT��\�������\��������Eԃ��Eԋ���������������\���;���������������;�����t6ha� ���wPh�`hL[�P�����h�`� ���wP������������;�����t
�  �  ��  �E����M�����,�����,����D;Dtǅ����   �
ǅ����    �������M��}� �  �E�����,���kU�kE�E��
��J�H�J�H�J�H�J�H�R�P�E�����,���kTU��Eԃ�k�M����B�A�B�A�B�A�B�A�R�Q�E�����,���kTU��Eԃ�k�M����B�A�B�A�B�A�B�A�R�Q�}� tB�E�����,���kTU��Eԃ�k�M����B�A�B�A�B�A�B�A�R�Q�E�����,���kU�kE�Eȋ
��J�H�J�H�J�H�J�H�R�P�E�����,����Uԉ�Eԃ��EԋE�����,���kTU�kE�Eȋ
��J�H�J�H�J�H�J�H�R�P�E�����,����UԉT�Eԃ��EԋE�����,���kTU�kE�Eȋ
��J�H�J�H�J�H�J�H�R�P�E�����,����UԉT�Eԃ��Eԃ}� t[�E�����,���kTU�kE�Eȋ
��J�H�J�H�J�H�J�H�R�P�E�����,����UԉT�Eԃ��E�� �E����M�����,�����,����D�D
�0����E�P蚞�����E�P莞�����n  �M�c���=  �[  �M�����������M�ҵ���������E�    �	�E����E��E�;�����}P�E��������<� u�ۋE��������|� t�E����������EԍP�M���E����������EԍLP��M�뜋�h�`� ��   PkM�Q����B���  �у�;��?����E��}� u3���  �E�PkM�Q�U�R�E�P��������h�`� ��   P��������Q����B���  �у�;������������������ u3��c  ������P��������Q������R������P��������Eԙ+���P�E�P�M葷����u"�E�P�������������P������3��  �M�n����EȋM�g���������ǅ����    ǅ����    �E�    �	�E����E��E�;������)  �E��������<� u��ǅ����    ������������������������M�������;���   ��������;E�}�������������T;U�|h�`� ��   P�$������   �����������k�M�k�����Uȋ��A�B�A�B�A�B�A�B�I�J���������������������������Tk�E�k�����Mȋ��P�Q�P�Q�P�Q�P�Q�@�A��������������������E��������|� ��   ��������;E�}�����������;E�|h�`� ��   P�1������   �����������k�M�k�����Uȋ��A�B�A�B�A�B�A�B�I�J��������������k�����E�k�����Mȋ��P�Q�P�Q�P�Q�P�Q�@�A���������������E�������������������������E�    �	�E����E��Eԙ+���9E�}#�E��������D�    �E���������   �Ǎ�����P�������E�P�������   �&�E�P��������E�P�������E�P������3�R��P�������XZ_^[��D  ;��E�����]Ë�   �����   G�����   A�����   4����   *�����   $�osadr pointsort ngonpointmap opadr sttpadr ��.�F�^���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �������Ef/Ev�E��Ef/Ev�E��E_^[��]�����������������������U����   SVW��@����0   �������EP���E�$�MQ�UR����HH���  �҃�;������_^[���   ;�������]��������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��a����E�     _^[���   ;��H�����]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;�������E�     _^[���   ;��������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��a����E�     _^[���   ;��H�����]��������������������������������������U����   SVW��@����0   �������EP����QH���  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��q����E�     _^[���   ;��X�����]��������������������������������������U����   SVW��@����0   �������EP����QH��  �Ѓ�;������_^[���   ;��������]������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;��h�����]��������������������������������������U����   SVW��@����0   �������E P�MQ���E�$�UR�EP�MQ����BH���   �у�;������_^[���   ;��������]���������������������������������U����   SVW��@����0   �������EP���E�$�MQ�UR�EP����QH���   �Ѓ�;��W���_^[���   ;��G�����]�������������������������������������U����   SVW��@����0   �������EP�MQ�UR����HH���  �҃�;������_^[���   ;��������]�����������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����BH���  �у�;��`���_^[���   ;��P�����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;������_^[���   ;��������]�������������������������U����   SVWQ������=   ������Y�M��E�    �E�    �E�    �E�8 u*�MQ�M�������uj�M��\�����uǅ���    �
ǅ���   �U�������E�8 uc�M������} u�EP�MQ�UR�EP�MQ�M�躖���7�E�E���M��}����E��}� t�EP�MQ�UR�E�P�MQ�M�胖���ыE�8 u�M��Y�����tǅ���    �
ǅ���   �M�������E�8 u�M��o����EP�M��Y����   �M��S����} u�EPj �MQ�UR�EP�M������E��uh  �#������E�}� u3��^�M�H���P�M��i����E�E���M�蘢���E��}� t1�EPj �MQ�U�R�EP�M�蠕���Eԃ}� t�E�P�M��W���뾋E�_^[���   ;��ʾ����]� �������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��`  �Ѓ�;������_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;�臽��_^[���   ;��w�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;�����_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;�苼��_^[���   ;��{�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��@_^[��]�����������������U����   SVWQ��4����3   ������Y�M���E�P����Q@�B,�Ѓ�;��^���_^[���   ;��N�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q@�B,�Ѓ�;�����_^[���   ;��޺����]����������������������������U����   SVWQ��0����4   ������Y�M���j�E�P����QH���   �Ѓ�;��y�����tǅ0���   �
ǅ0���    ��0���_^[���   ;��I�����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��!��E��HQ����Bl�H�у�;��ι��_^[���   ;�边����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;��[���_^[���   ;��K�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M��QR����Hl�Q�҃�;��ܸ��_^[���   ;��̸����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;��[���_^[���   ;��K�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��  �҃�;�����_^[���   ;��Է����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��  �҃�;��d���_^[���   ;��T�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���j �E�P����QH���   �Ѓ�;�����_^[���   ;��ٶ����]�����������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;��{���_^[���   ;��k�����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��T  �Ѓ�;�����_^[���   ;��������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��  �у�;�藵��_^[���   ;�臵����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����HH���  �҃�;�����_^[���   ;��������]� �����������������������������������U����   SVWQ��0����4   ������Y�M��E��x ~�   k� �U�
芄����0����
ǅ0���������0���_^[���   ;��i�����]���������������������������������������U����   SVWQ��(����6   ������Y�M�j h�  �M��W~�����T����E�M�褡�����}�u�E���3�_^[���   ;��׳����]�������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��(  �Ѓ�;��k���_^[���   ;��[�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP���E�$�MQ�U�R����HH��0  �҃�;�����_^[���   ;��ײ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M����   ��;��g���_^[���   ;��W�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QH���  �Ѓ�;��߱��_^[���   ;��ϱ����]� ��������������������������U����   SVWQ������9   ������Y�M��E�P�M�Q�UR�EP�M�迧���E�;Eu�E����E�;Eu�E�����R��P��������XZ_^[���   ;��4�����]� �I    ������   �����   �l2 l1 ������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��  �Ѓ�;�苰��_^[���   ;��{�����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��8  �у�;�觯��_^[���   ;�藯����]� ����������������������������������U����   SVWQ������;   ������Y�M���E�P�����Q����BH��\  �у�;��$����U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;�������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;��w���_^[���   ;��g�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;������_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M�h�  �M�����_^[���   ;�菭����]�����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;��+���_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;�軬��_^[���   ;�諬����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M��QR����Hl�Q�҃�;��H���_^[���   ;��8�����]� �����������������������������������U����   SVWQ��4����3   ������Y�M�h�  �M��\���_^[���   ;��ϫ����]�����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��  �Ѓ�;��k���_^[���   ;��[�����]�������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M��{���_^[���   ;��������]���������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��  �Ѓ�;�蛪��_^[���   ;�苪����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���  �҃�;��$���_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��P  �Ѓ�;�諩��_^[���   ;�蛩����]�������������������������U����   SVWQ��4����3   ������Y�M�����E�$�EP����Q�M����   ��;��.���_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��4  �Ѓ�;�軨��_^[���   ;�諨����]�������������������������U����   SVWQ��4����3   ������Y�M���j�E�P����QH���   �Ѓ�;��I���_^[���   ;��9�����]�����������������������U����   SVWQ��4����3   ������Y�M�h(  �M��l���_^[���   ;��ߧ����]�����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��,  �҃�;��t���_^[���   ;��d�����]� �������������������������������U����   SVWQ��4����3   ������Y�M�j h(  �M��(���_^[���   ;��������]���������������������������U���,  SVWQ�������K   ������Y�M���t���E�}� t�} u3���   �M��2|���E��M�舻�����Eԃ}� u�E���   �E�    �	�Eȃ��EȋM�����9E���   �E�P�M�Q�U�R�E�P�M�]�����u�ȋE��E��	�E����E��E�;E�_�E�����u$�E������M������U��u��D;Du���E���P�M�Of���M����T��U��}��t�E�P�M��bk����K����E�R��P����U���XZ_^[��,  ;�蘥����]� �I    ������   ������   ��b a ������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�    �}u�M�萸���E��$�} u�M��T����E���}u�M������E�}� u3���E�P�MQ�M��}��_^[���   ;��t�����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��  �у�;������_^[���   ;�������]� ����������������������������������U����   SVWQ������;   ������Y�M���EP�MQ���E�$�U�R�����P����QH��  �Ѓ�;��_����M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;��'�����]� ��������������������������������������������������U����   SVWQ������;   ������Y�M���EP�MQ���E�$�U�R�����P����QH��  �Ѓ�;�菢���M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;��W�����]� ��������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��\  �Ѓ�;��ۡ��_^[���   ;��ˡ����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���   �҃�;��d���_^[���   ;��T�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;�����_^[���   ;��נ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��p  �҃�;��d���_^[���   ;��T�����]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��  �҃�;�����_^[���   ;��ԟ����]� �������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��B��;��p���_^[���   ;��`�����]������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;������_^[���   ;�������]�������������������������U����   SVWQ������;   ������Y�M���EP�MQ�����R����P�M����   ��;�聞���M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[���   ;��I�����]� ������������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����QH���   �Ѓ�;��ȝ��_^[���   ;�踝����]��������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P����QH�B�Ѓ�;��A���_^[���   ;��1�����]� ����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��X  �Ѓ�;��˜��_^[���   ;�軜����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��,  �Ѓ�;��[���_^[���   ;��K�����]�������������������������U����   SVWQ��4����3   ������Y�M��E���U����k��_^[���   ;�������]� �����������������������U����   SVWQ��4����3   ������Y�M��E�� %�����_^[��]��������������������������U����   SVWQ��0����4   ������Y�M���E��HQ����Bl�H�у�;��;����} u�   �T��EP�MQ�UR�EP����Ql��Ѓ�;������M��A�E��x tǅ0���   �
ǅ0���    ��0���_^[���   ;��ʚ����]� �����������������������������������������������������U����   SVWQ��0����4   ������Y�M���EP����QH��x  �Ѓ�;��K����M���E��8 tǅ0���   �
ǅ0���    ��0���_^[���   ;�������]� ���������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QH��   �Ѓ�;�菙��_^[���   ;�������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���   �҃�;�����_^[���   ;�������]� �������������������������������U����   SVW��@����0   �������E0P�M,Q�U(R�E$P�M Q���E�$���E�$�UR�EP����QH��P  �Ѓ�,;��n���_^[���   ;��^�����]��������������������������������������������U����   SVWQ��4����3   ������Y�M�j h�  �M��$������h��_^[���   ;�������]��������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;�臗��_^[���   ;��w�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E���U���vt��_^[���   ;�������]� �����������������������U����   SVWQ��0����4   ������Y�M��E����   �uǅ0���   �
ǅ0���    ��0���_^[��]������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H,�у�;��:���_^[���   ;��*�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH���   �҃�;�贕��_^[���   ;�褕����]� �������������������������������U����   SVW��@����0   ������E;E}�E��E;E~�E��E_^[��]�������������������������������U����   SVWQ��(����6   ������Y�M��EP�s�����E�}� t�EP�M�Q�M��PX���E�_^[���   ;��Ĕ����]� �������������������������������U����   SVWQ��(����6   ������Y�M��EP�MQ��t�����E�}� t�EP�M�Q�M���W���E�_^[���   ;��@�����]� ���������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;��ۓ��_^[���   ;��˓����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��t  �Ѓ�;��k���_^[���   ;��[�����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��   �҃�;������_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;��w���_^[���   ;��g�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��  �҃�;������_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QH��   �Ѓ�;��o���_^[���   ;��_�����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����BH��|  �у�;�����_^[���   ;��ې����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HH��8  �҃�;��d���_^[���   ;��T�����]� �������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P����QH��t  �Ѓ�;��ޏ��_^[���   ;��Ώ����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;��g���_^[���   ;��W�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H@�Q(�҃�;�����_^[���   ;��׎����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���  �Ѓ�;��k���_^[���   ;��[�����]�������������������������U����   SVWQ��4����3   ������Y�M���EPj�M�Q����BH���   �у�;������_^[���   ;�������]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EPj �M�Q����BH���   �у�;��u���_^[���   ;��e�����]� ��������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P����QH��h  �Ѓ�;�����_^[���   ;��ތ����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���   �у�;��w���_^[���   ;��g�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��B|��;������_^[���   ;�������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��p  �у�;�臋��_^[���   ;��w�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;�����_^[���   ;��������]� ����������������������������������U���   SVWQ�� ����@   ������Y�M�j h�  �M��ba���} u�   �uj h�  �M��xW���E�}� u3��Y�M��L���EPh�  �M���V�����E�$h�  �M�聚��j �E�P�M��V��ǅ���   �M��qN�������R��P�,�距��XZ_^[��   ;��������]� �   4�����   @�bc �������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��X  �у�;��W���_^[���   ;��G�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��d  �у�;��׈��_^[���   ;��ǈ����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EPj�M�Q����BH���   �у�;��U���_^[���   ;��E�����]� ��������������������������������U����   SVWQ������?   ������Y�M��M��]���E�}� u3��j  �E�    �}u�M�蘛���E��$�} u�M��\t���E���}u�M�������E��}� u3��  �M�蔘���E�    �	�Eԃ��EԋM��q���9E���   �E�P�M��G���Eȃ}� u�ϸ   k� �UȋD
P�M�*o����t�E���P�M���L���   �� �MȋTR�M��n����t�Eԍ�   Q�M��L���E����M����U�u�D;Dt.�   ���MȋTR�M�n����t�Eԍ�   Q�M��RL���   k��UȋD
P�M�n����t�Eԍ�   Q�M��#L��������   _^[���   ;��j�����]� ���������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;�觅��_^[���   ;�藅����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��PH��;��*���_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P����QH��l  �Ѓ�;�螄��_^[���   ;�莄����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����BH���  �у�;�����_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�UR�E�P����QH���  �Ѓ�;�胃��_^[���   ;��s�����]� ������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;�����_^[���   ;��������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;�蛂��_^[���   ;�苂����]�������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����QH���  �Ѓ�;��$���_^[���   ;�������]����������������������������������U����   SVWQ��4����3   ������Y�M���EP���E�$�M�Q����BH���  �у�;�蚁��_^[���   ;�芁����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R����HH���  �҃�0;������_^[���   ;��������]�, �������������������������������������������U����   SVW��@����0   �������E0P���E(�$�M$Q�U R�EP�MQ�UR�EP�MQ�UR����HH���  �҃�,;��D���_^[���   ;��4�����]����������������������������������U����   SVWQ��4����3   ������Y�M���E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R����HH���  �҃�0;����_^[���   ;������]�, �������������������������������������������U����   SVW��@����0   �������E P�MQ�UR�EP�MQ�UR�EP����QH���  �Ѓ�;����_^[���   ;���~����]��������������������������������������U����   SVWQ��4����3   ������Y�M�����E�$�E�P����QH��$  �Ѓ�;��~~��_^[���   ;��n~����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��H  �у�;��~��_^[���   ;���}����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��L  �Ѓ�;��}��_^[���   ;��{}����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��<  �у�;��}��_^[���   ;��}����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����QH��@  �Ѓ�;��|��_^[���   ;��|����]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH���  �у�;��|��_^[���   ;��|����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��  �у�;��{��_^[���   ;��{����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH��T  �Ѓ�;��{��_^[���   ;��{����]�������������������������U����   SVWQ��4����3   ������Y�M��?���M���E�_^[���   ;��z����]�����������������������������U����   SVWQ��4����3   ������Y�M��E�P�r>�����E��     _^[���   ;��Gz����]���������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]������������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]�����������̋�`��`��`��`��`��`��` ��`��������������U����   SVWQ��0����4   ������Y�M��M�������tǅ0���   �
ǅ0���    ��0���_^[���   ;��$y����]����������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��M��}���E_^[���   ;��x����]� ����������������������������U����   SVWQ��4����3   ������Y�M��   @_^[��]� ���������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U���  SVW��x����b   ������} u3��   j h�   ��<���P�;O�����E��\����E��|����E�E��E��<���ǅ@���d�E�)8�E�%P�E��T�E��M�E��T�E��M�E��8�E��bh�   ��<���P�MQ�URj�E����R��P��������XZ_^[�Ĉ  ;��<v����]Ð   ��<����   ��np �����������������������������������������������������������������U����  SVW��(����v   ������ǅ ���    �}( uǅ0���    �M�]����0����!  �E�    �M��~������  �M���I���M��5?������   �EP��H�����_���� ���j h|`�������kQ���� ���P��l����_���� ���j j���H���Q��l���R������P��`������ ���P������Q�n������ ���P������R�n������ ��� P�M��7������6����uǅ(���   �
ǅ(���    ��(�����?����� ����� t�� ���ߍ�������;���� �����t�� ��������;���� �����t�� �����������;���� �����t�� ������l����~;���� �����t�� �����������\���� �����t�� ������H����D;����?�����t(�E(P�M$Q�M��=��P�UR�EP�MQ��Y�����E��M��H~���!�E(P�M$Qj �UR�EP�MQ�Y�����E��E�������M�[�������R��P�������XZ_^[���  ;��Rs����]ÍI    ������   ��icon �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���  SVW��x����b   ������j h�   ��<���P�J����ǅ\���    �E��|���h�   ��<���P�MQ�URj�]A����R��P�,�超��XZ_^[�Ĉ  ;���q����]Ë�   4�<����   @�np ���������������������������������������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVW��@����0   ������E������� _^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��E��M���j j j �E��Q����B�H�у�;���p���U��B�E�_^[���   ;��p����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H|�Q�҃�;��Gp��_^[���   ;��7p����]� ����������������������������������U����   SVWQ��(����6   ������Y�M���E�P������   �BX�Ѓ�;���o���E�}� u3���EP�MQ�M��m��_^[���   ;��o����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H|�Q8�҃�;��'o��_^[���   ;��o����]� ����������������������������������U����   SVWQ��(����6   ������Y�M���E�P������   �BX�Ѓ�;��n���E�}� u3���EP�MQ�M��I��_^[���   ;��~n����]� �����������������������������������������U����   SVWQ��4����3   ������Y�M��E��x u3��9��E��HQ�UR�EP�M��R����H�Q�҃�;���m���M��A�   _^[���   ;���m����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���j j j �E��Q����B�H�у�;��fm���U��B_^[���   ;��Pm����]������������������������������U����   SVWQ��(����6   ������Y�M�j\�  ���E�}� t	�E�x\ u�<��E�P�M�Q\�҃�;���l���EP�M��4]���EP�M���2���EP�M���2���E�_^[���   ;��l����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�j\��  ���E�}� t	�E�x\ u�0��E�P�M�Q\�҃�;��l���EP�M��t\���EP�M��2���E�_^[���   ;���k����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j\�F  ���E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;��fk���EP�M���[���E�_^[���   ;��Gk����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�j\�  ���E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;���j���EP�M��=L���E�_^[���   ;��j����]� ����������������������������������U����   SVWQ������;   ������Y�M�j\�  ���E�}� t	�E�x\ u�0��E�P�M�Q\�҃�;��&j���EP������[��P�M��xZ���E�_^[���   ;���i����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j\�V  ���E�}� t	�E�x\ u���E�P�M�Q\�҃�;��vi���E�_^[���   ;��ci����]���������������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]��������������������U����   SVWQ��(����6   ������Y�M�j`�  ���E�}� t	�E�x` u���E�P�M�Q`�҃�;��h��_^[���   ;��h����]������������������������������������U����   SVWQ��(����6   ������Y�M�jx��  ���E�}� t	�E�xx u�E����E�P�MQ�U�Bx�Ѓ�;��h���E�_^[���   ;���g����]� ���������������������������������������U����   SVWQ������:   ������Y�M�jt�V  ���E�}� t	�E�xt uh���M��Z���E�:��EP�M�Q�����R�E�Ht�у�;��[g��P�M�T���������d���E_^[���   ;��4g����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�j|�
  ���E�}� t	�E�x| u3����E�P�MQ�U�B|�Ѓ�;��f��_^[���   ;��f����]� �������������������������������������������U����   SVWQ��0����4   ������Y�M��E�M��;t3���   �E�x uN�E�8 uF�E�x u=�E��x u�M��9 u�U��z uǅ0���   �
ǅ0���    ��0����   �R�E��x uI�E��8 uA�E��x u8�E�x u�M�9 u�U�z uǅ0���   �
ǅ0���    ��0����M�E�x t�E��x t�E�M��P;Qt3��)�E�x t�E��x t�E�M��P;Qt3���   _^[��]� �������������������������������������������������������������������������������������������U����   SVWQ��$����7   ������Y�M�j|�V  ���E�}� t	�E�x| u�   �<��E�P�MQ�U�B|�Ѓ�;��md����uǅ$���   �
ǅ$���    ��$���_^[���   ;��=d����]� ����������������������������������������U����   SVWQ��0����4   ������Y�M��EP�M���x����uǅ0���   �
ǅ0���    ��0���_^[���   ;��c����]� ���������������������������U����   SVWQ��(����6   ������Y�M�jp�  ���E�}� t	�E�xp u������EP�M�Q�U�Bp�Ѓ�;��-c��_^[���   ;��c����]� ����������������������������������������U����   SVW��$����7   ������h�   �x  ���E��}� t�E����    u�EP�M��O���E�=��EP�MQ��(���R�E����   �у�;��xb��P�M�O����(�����_���E_^[���   ;��Qb����]�����������������������������������������������U����   SVWQ������:   ������Y�M�h�   �  ���E�}� t�E샸�    u�E��4��EP�M�Q�����R�E싈�   �у�;��a��������._���E�_^[���   ;��a����]� ��������������������������������������������U����   SVW��4����3   ������j��  ���E��}� t	�E��x u3���E���H��;��a��_^[���   ;�� a����]������������������������������U����   SVWQ������?   ������Y�M�h�   �c  ���E�}� t�E샸�    uj ������R��P�M��S���E�9��EP�����Q�U�M����   ��;��]`��P�M�M���������]���E_^[���   ;��6`����]� �������������������������������������������������U����   SVWQ��(����6   ������Y�M�j<�  ���E�}� t	�E�x< u���EP�M�Q�U�B<�Ѓ�;��_��_^[���   ;��_����]� �����������������������������U����   SVWQ��(����6   ������Y�M�h�   ��  ���E�}� t�E샸�    u���EP�U�M����   ��;��_��_^[���   ;���^����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S  ���E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��c^��_^[���   ;��S^����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�j4�  ���E�}� t	�E�x4 u3����E�P�M�Q4�҃�;���]��_^[���   ;��]����]����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �  ���E�}� t�E샸�    u3����E�M����   ��;��/]��_^[���   ;��]����]���������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �s   ���E�}� u3��'��EP�MQ�UR�E�P�M싑�   �҃�;��\��_^[���   ;��{\����]� ��������������������������������������U����   SVW��@����0   ������h���EPhD ��A����_^[���   ;��\����]�������������������������U����   SVWQ��(����6   ������Y�M�h�   �s������E�}� t�E샸�    u3����EP�U�M����   ��;��[��_^[���   ;��{[����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�jD��������E�}� t	�E�xD u3����E�P�M�QD�҃�;���Z��_^[���   ;���Z����]����������������������������������U����   SVWQ��(����6   ������Y�M�jL�F������E�}� u3����EP�M�Q�U�BL�Ѓ�;��iZ��_^[���   ;��YZ����]� ������������������������������������U����   SVW������9   ������h�   �������E��}� u�M�_���E�9��EP�� ���Q�U����   �Ѓ�;���Y��P�M�P6���� �����A���E_^[���   ;��Y����]���������������������������������������������������U����   SVW��4����3   ������j��������E��}� t	�E��x u3�� ��EP�MQ�UR�E��H�у�;��Y��_^[���   ;��Y����]�������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;��sX��_^[���   ;��cX����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�U�M����   ��;���W��_^[���   ;��W����]� ��������������������������������������U����   SVW��4����3   ������E�8 u�?j�������E��}� t	�E��x u�!��EP�M��Q�҃�;��1W���E�     _^[���   ;��W����]��������������������������������������U����   SVWQ��(����6   ������Y�M�jH�v������E�}� u���EP�M�Q�U�BH�Ѓ�;��V��_^[���   ;��V����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M��E�    �	�E���E�E�P�M��Y*���8 t��E�_^[���   ;��V����]����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� u�'��EP�MQ�UR�E�P�M싑�   �҃�;��}U��_^[���   ;��mU����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�j$��������E�}� t	�E�x$ u3����E�P�M�Q$�҃�;���T��_^[���   ;���T����]����������������������������������U����   SVWQ������9   ������Y�M�h�   �3������E�}� t�E샸�    u3����E�M����   ��;��OT���E��E�_^[���   ;��9T����]���������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� u3����EP�M�Q�U싂�   �Ѓ�;��S��_^[���   ;��S����]� ������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� u3����EP�M�Q�U싂�   �Ѓ�;��#S��_^[���   ;��S����]� ������������������������������U����   SVWQ��(����6   ������Y�M�j8�v������E�}� t	�E�x8 u3��(��EP�MQ�UR�EP�M�Q�U�B8�Ѓ�;��R��_^[���   ;��tR����]� �����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� u3����EP�M�Q�U싂�   �Ѓ�;���Q��_^[���   ;���Q����]� ������������������������������U����   SVWQ��(����6   ������Y�M�j(�6������E�}� t	�E�x( u3��$��EP�MQ�UR�E�P�M�Q(�҃�;��HQ��_^[���   ;��8Q����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�j,�������E�}� t	�E�x, u3�� ��EP�MQ�U�R�E�H,�у�;��P��_^[���   ;��P����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�jP��������E�}� u3�� ��EP�MQ�U�R�E�HP�у�;��P��_^[���   ;��P����]� ��������������������������������U����   SVWQ��(����6   ������Y�M�jT�f������E�}� u3����E�P�M�QT�҃�;��O��_^[���   ;��}O����]���������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� u3��/��EP�MQ�UR�EP�MQ�U�R�E싈�   �у�;���N��_^[���   ;���N����]� ����������������������������������������������U����   SVWQ��$����7   ������Y�M��E�    �	�E���E�E�P�M��"���8 t(�E�P�M�"��P�M�Q�M��"�����[����t�뾃} t�E�M��}� ~�E�P�M��\"���8 uǅ$���   �
ǅ$���    ��$���_^[���   ;���M����]� �����������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j�6������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;��PM��_^[���   ;��@M����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�M�Q�U�B�Ѓ�;��L��_^[���   ;��L����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M��} u3��@j��������E�}� t	�E�x u3�� ��EP�MQ�U�R�E�H�у�;��L��_^[���   ;���K����]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�jl�F������E�}� t	�E�xl u���E�P�M�Ql�҃�;��fK��_^[���   ;��VK����]������������������������������������U����   SVWQ��(����6   ������Y�M�jh�������E�}� t	�E�xh u���EP�M�Q�U�Bh�Ѓ�;���J��_^[���   ;���J����]� �����������������������������U����   SVWQ��(����6   ������Y�M�h�   �#������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;��7J��_^[���   ;��'J����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3����EP�U�M����   ��;��I��_^[���   ;��I����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;���H��_^[���   ;���H����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�jd�6������E�}� t	�E�xd u���EP�M�Q�U�Bd�Ѓ�;��RH��_^[���   ;��BH����]� �����������������������������U����   SVWQ��(����6   ������Y�M�j(�������E�}� t	�E�x0 u3��$��EP�MQ�UR�E�P�M�Q0�҃�;��G��_^[���   ;��G����]� �����������������������������������U����   SVWQ��(����6   ������Y�M�jX�������E�}� u���EP�M�Q�U�BX�Ѓ�;��+G��_^[���   ;��G����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�j �v������E�}� t	�E�x  u3����E�P�M�Q �҃�;��F��_^[���   ;��F����]����������������������������������U����   SVWQ��(����6   ������Y�M�h�   ��������E�}� t�E샸�    u3����EP�M�Q�U싂�   �Ѓ�;���E��_^[���   ;���E����]� ����������������������������������U����   SVW��<����1   ������E��<�����<���t��E����E����   _^[��]� ��������������������������������U����   SVW������:   ������E�����������������������q  ������$���   �]  ���������=����   �EP�E����=�2  }
������&  �} u
������  h@a�$���Ph��j������� ����� ��� t�� ����t��������
ǅ���    ���������=�� t�EP����<!���   �   �EP�MQ��J������u����   �   �|�D���u��������u\�X0���@���=�� t?�����8�����8�����,�����,��� tj��,����:��������
ǅ���    ���    �   ����_^[���   ;��C����]Ð* ������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��M������E�    �	�E���E�}�}�E�M��D�    ��E�_^[���   ;��B����]���������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �M��A    �U��B    �E��@    �E��@    �E�_^[��]�����������������������������������������U����   SVWQ��4����3   ������Y�M��M����R;���M��qF���E�_^[���   ;��A����]��������������������U����   SVWQ��4����3   ������Y�M��M����_^[���   ;��4A����]������������������U����   SVWQ��4����3   ������Y�M��M�����M����'��_^[���   ;���@����]�����������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B��(  �у�;��w@���E�_^[���   ;��d@����]� �������������������������������U����   SVWQ��4����3   ������Y�M���E�P�MQ����B��,  �у�;���?��_^[���   ;���?����]� ����������������������������������U����   SVWQ��0����4   ������Y�M���E�P�MQ����B��,  �у�;��w?����uǅ0���   �
ǅ0���    ��0���_^[���   ;��G?����]� ����������������������������������U����   SVW��@����0   ������E#E_^[��]����������������������U����   SVWQ��4����3   ������Y�M��M���S���E��t�E�P�qR�����E�_^[���   ;��>����]� ������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H�Q@�҃�;��'>��_^[���   ;��>����]� ����������������������������������U����   SVW��@����0   �����󫡸��H����;��=��_^[���   ;��=����]��������������������������U����   SVW��@����0   �����󫡸��H���   ��;��X=��_^[���   ;��H=����]����������������������U����   SVW��@����0   �����󫡸��H��   ��;���<��_^[���   ;���<����]����������������������U����   SVW��@����0   �����󫡸��H��\  ��;��<��_^[���   ;��<����]����������������������U����   SVW��0����4   ������h�a�(���Ph��h�   �O������8�����8��� t��8����tH����0����
ǅ0���    ��0���_^[���   ;���;����]���������������������������������������������U����   SVW��@����0   �����󫡸��H����;��;��_^[���   ;��|;����]��������������������������U����   SVWQ��4����3   ������Y�M��EP�M��P��_^[���   ;�� ;����]� ���������������������������U����   SVWQ��4����3   ������Y�M��EP�M��O��_^[���   ;���:����]� ���������������������������U����   SVWQ��4����3   ������Y�M��M�������xX u�'��EP�M���������M�������H �WX��;��E:��_^[���   ;��5:����]� ��������������������������������U����   SVWQ��4����3   ������Y�M���EP�M��N������M��D����H �WH��;���9��_^[���   ;��9����]� ��������������������������������U����   SVWQ��4����3   ������Y�M��M�������xT u����+��EP�MQ�M��������M������H �WT��;��.9��_^[���   ;��9����]� �����������������������������������������U���  SVWQ�������C   ������Y�M��} t<�M�������E�P�M�� ������M������H �WL��;��8���M��M�������} t?�������<>��P�M�$���������} ���M�������@@�EЃ}� t�E�P�M��#��R��P�(��K��XZ_^[��  ;��$8����]� �I    (����   (bc ���������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M������xL u3��/��EP�MQ�UR�M���������M�������H �GL��;��[7��_^[���   ;��K7����]� ��������������������������������������U����   SVWQ��4����3   ������Y�M��M��d����x` u� }  �'��EP�M��I������M��?����H �W`��;���6��_^[���   ;��6����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��M�������xH u3��#�M��������M��������H �FH��;��'6��_^[���   ;��6����]�������������������������������������U����   SVWQ��4����3   ������Y�M��M��4����xX u����'��EP�M��������M������H �WX��;��5��_^[���   ;��5����]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��������M������H �G@��;��5��_^[���   ;���4����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M��������M�������H �GD��;��}4��_^[���   ;��m4����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��M������xP u����3��EP�MQ�UR�EP�M��_������M��U����H �WP��;���3��_^[���   ;���3����]� ���������������������������������U����   SVWQ��4����3   ������Y�M��M�������xP u������;��EP�MQ�UR�EP�MQ�UR�M��������M������H �GP��;��,3��_^[���   ;��3����]� ���������������������������������������U����   SVWQ��$����7   ������Y�M�j�EP��<������tǅ$���   �
ǅ$���    ��$���Q�M��-���E�M����;E��M�J=��;E�~������3��EP�MQ�UR�EP�M���������M������H �WD��;��>2��_^[���   ;��.2����]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��4����xT u������+��EP�MQ�M��������M������H �WT��;��1��_^[���   ;��|1����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��l  �у�;��1��_^[���   ;���0����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H�Q�҃�;��0��_^[���   ;��w0����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�M���:����P�M��P����Pj j �E�P����Q�B4�Ѓ� ;���/��_^[���   ;���/����]� ���������������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q����B�H4�у� ;��R/��_^[���   ;��B/����]� �����������������������������U����   SVWQ��4����3   ������Y�M��M������M���3��_^[���   ;���.����]��������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��~.��_^[���   ;��n.����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H��h  �҃�;���-��_^[���   ;���-����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H���   �҃�;��h-��_^[���   ;��X-����]� �����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�H\�у�;���,��_^[���   ;���,����]� �������������������������������������U����   SVWQ��0����4   ������Y�M��} t�M�D�����0����
ǅ0���    ��0���P�M�Q����B��8  �у�;��D,��_^[���   ;��4,����]� �����������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B �Ѓ�;��+��_^[���   ;��+����]����������������������������U����   SVWQ��4����3   ������Y�M��M��S���_^[���   ;��T+����]������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;��+����]������������������U����   SVW��@����0   �������E�Q����B�H�у�;��*���E�     _^[���   ;��*����]��������������������������������������U����   SVW��@����0   �������E�Q����B���   �у�;��.*���E�     _^[���   ;��*����]�����������������������������������U����   SVW��@����0   �������E�Q����B��$  �у�;��)���E�     _^[���   ;��)����]�����������������������������������U����   SVW��@����0   �������E�Q����B��`  �у�;��.)���E�     _^[���   ;��)����]�����������������������������������U����   SVW��$����7   ������E�8 t?�E���8�����8�����,�����,��� tj��,��������$����
ǅ$���    �E�     _^[���   ;��q(����]�����������������������������������������������U����   SVW��@����0   �������E�Q����B�H�у�;��(���E�     _^[���   ;���'����]��������������������������������������U����   SVW��@����0   �������E�Q����B�H�у�;��'���E�     _^[���   ;��h'����]��������������������������������������U����   SVWQ��4����3   ������Y�M��E��8 t j j j�E���P�M��	�K���E��     �E��x` t�E���`P�������_^[���   ;���&����]������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q���   �Ѓ�;��[&��_^[���   ;��K&����]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;���%��_^[���   ;���%����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��~%��_^[���   ;��n%����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�BP�Ѓ�;��%��_^[���   ;���$����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�HT�у�;��$��_^[���   ;��$����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�HT�у�;��$��_^[���   ;��
$����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�B�Ѓ�;��#��_^[���   ;��#����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B�HX�у�;��#��_^[���   ;��#����]� �������������������������U����   SVWQ������<   ������Y�M���h�  �E�P�� ���Q����B���   �у�;��"�����]��������� ����Z��������_^[���   ;��q"����]�����������������������������������������������U����   SVWQ������9   ������Y�M���EP�MQ�U�R�� ���P����Q���   �Ѓ�;���!��P�M������ ��������E_^[���   ;���!����]� ��������������������������������U����   SVW��@����0   �����󫡸��H��t  ��;��h!��_^[���   ;��X!����]����������������������U����   SVW��@����0   �����󫡸��H��4  ��;��!��_^[���   ;��� ����]����������������������U����   SVW��@����0   �����󫡸��H��p  ��;�� ��_^[���   ;�� ����]����������������������U����   SVW��@����0   �����󫡸��H��0  ��;��H ��_^[���   ;��8 ����]����������������������U����   SVWQ������9   ������Y�M���EP�M�Q�� ���R����H��L  �҃�;�����P�M�U����� ��������E_^[���   ;������]� �������������������������������������U����   SVWQ��4����3   ������Y�M��} t�E�M��Ap� �E��xd t�E��@h��E��x|u�   �3�_^[��]� ����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�BL�Ѓ�;����_^[���   ;������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�BL�Ѓ�;��N��_^[���   ;��>����]����������������������������U����   SVWQ������<   ������Y�M��M�S-���M�������uh�a�0���P�_/����3��   �E�    ��E�P�M�Q�UR�E�P����Q���   �Ѓ�;������u3��M�E�    �	�Eԃ��EԋE�;E�}"�EԋM��<� u��EԋM���R�M�&���͍E�P��������   R��P�C��0��XZ_^[���   ;��!����]�    C����   (C����   $Carr count ����������������������������������������������������������������������������������U����   SVWQ������<   ������Y�M��M�	����M��.�����uh�a�4���P��-����3��   �E�    ��E�P�M�Q�UR�E�P����Q���   �Ѓ�;������u3��i�}� u3��_�E�    �	�Eԃ��EԋE�;E�}4�EԋM��<� t�EԋM���������u�ϋEԋM���R�M�8���뻍E�P�'������   R��P��D�B/��XZ_^[���   ;������]�    �D����   �D����   �Darr count ��������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M�����P��M���|  ��;�����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q��T  �Ѓ�;��K��_^[���   ;��;����]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q�B�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B���   �у�;��K��_^[���   ;��;����]� ��������������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQ����B��   �у�;�����_^[���   ;������]������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@`    �E��@d    �E��@h    �E��x^�@p�E��@x�����E��@|   _^[��]��������������������������������������������U����   SVW�� ����8   ������M������E�P�MQ�i$������t�}� u3���E�P�M�Q�U�R�E�P�M������R��P��H�/+��XZ_^[���   ;��r����]ÍI    �H����   �Hdat ����������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q��P  �Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q�Bh�Ѓ�;��n��_^[���   ;��^����]����������������������������U����   SVWQ��4����3   ������Y�M��E��8 th�a�,���P�'�����E��x` th�a�,���P�l'�����M��c����M�����E�P�M���dQ�U��BxP�MQ�U���`R��������M��A|�E��x|u�E��8 u>�E��8 u�E��x|u
�E��@|�����E��     �E���`P�r������E��@|�   �E��xd ��   �E���pP�M���hQ�UR�t������u0�E��@h    �E��x^�@ph�a�,���P�&�����EP�M��������j j j�E���P�M��	�"����U��B|�E��x|t�M��I����E��@|��E��@x�����E��@|_^[���   ;������]� ����������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���E P�MQ�UR�EP�MQ�UR�EP�M�Q����B�H�у� ;�����_^[���   ;������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��<  �у�;��G��_^[���   ;��7����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q��@  �Ѓ�;����_^[���   ;������]� ��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ�U�R����H��d  �҃�;��8��_^[���   ;��(����]� �����������������������������������U����   SVWQ��4����3   ������Y�M��E��xd u�E��@`�}�E��M;Hxu�E��@`�j�EP�M��Q`Rj�E���P�M��	������U��B|�E��x|u �E��M�Hx�} t	�E�    �E��@`��E��@x�����} t�E�M��Q|�3�_^[���   ;��>����]� ���������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�HD�у�;����_^[���   ;������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q�M��B$��;��2��_^[���   ;��"����]� �����������������������������U����   SVWQ��4����3   ������Y�M���E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P����Q�B`�Ѓ�(;����_^[���   ;������]�$ �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B�H,�у�;����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B���   �у�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B�H(�у�;����_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H���   �҃�;����_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��X  �у�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M���x  ��;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B�H�у�;����_^[���   ;��
����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B��H  �у�;����_^[���   ;������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H��D  �҃�;����_^[���   ;������]� �������������������������������U����   SVWQ��4����3   ������Y�M��E��@    �E��     �E��@    �E��@   �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP����Q@�M����   ��;��
��_^[���   ;��
����]� ��������������������������U����   SVW��@����0   �����󫡸��H|��Q ��;��	��_^[���   ;��	����]�������������������������U����   SVW��@����0   �����󫡸��H|����;��\	��_^[���   ;��L	����]��������������������������U����   SVW��@����0   �������EP����Q@���   �Ѓ�;�����_^[���   ;�������]������������������������������U����   SVW��@����0   �����󫡸��H@��Q0��;����_^[���   ;��{����]�������������������������U����   SVW��@����0   �����󫡸��H@��Q0��;��+��_^[���   ;������]�������������������������U����   SVW��@����0   �������j�EPj ����Q@�B4�Ѓ�;����_^[���   ;������]�����������������������������U����   SVW��@����0   �������EP�MQj ����B@�H4�у�;��M��_^[���   ;��=����]���������������������������U����   SVW��@����0   �������j�EPh   @����Q@�B4�Ѓ�;�����_^[���   ;�������]��������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M����   ��;��k��_^[���   ;��[����]� ����������������������U����   SVW��@����0   ������h��hE  �M�6������������Ph��hE  �M����������P����H��T  �҃�;�����_^[���   ;�������]�����������������������������������������������U����   SVW��@����0   �������EP�MQ����B��T  �у�;��L��_^[���   ;��<����]��������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ������   �M����   ��;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M��BT��;��c��_^[���   ;��S����]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��B|��;��~��_^[���   ;��n����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P@�M����   ��;����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��BX��;����_^[���   ;��~����]� �������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B|�H(�у�;�����E�     _^[���   ;�� ����]������������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B|�H�у�;�����E�     _^[���   ;������]������������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B@�H�у�;�����E�     _^[���   ;�� ����]������������������������������U����   SVW��@����0   ������E�8 t ��E�Q����B@�H�у�;�� ���E�     _^[���   ;�� ����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�MQ������   �M����   ��;�� ��_^[���   ;��������]� �����������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M��Bt��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q@�BH�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M����   ��;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ������   �M��P��;��'���_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��B$��;�����_^[���   ;�������]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP������   �M����   ��;��,���_^[���   ;�������]� ���������������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M��Bx��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BH��d  �у�;��7���_^[���   ;��'�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QH���   �Ѓ�;�����_^[���   ;�������]�������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M��Pl��;��J���_^[���   ;��:�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��Bd��;������_^[���   ;�������]� �������������������������U����   SVWQ��4����3   ������Y�M�������   ��M��Bt��;��`���_^[���   ;��P�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M����   ��;������_^[���   ;��������]� �����������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M����   ��;��p���_^[���   ;��`�����]������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M��B��;������_^[���   ;��������]� �������������������������������U����   SVWQ��4����3   ������Y�M�����P@��M����   ��;�����_^[���   ;��p�����]������������������������������U����   SVW��4����3   ������}qF t�1�E�E��}� u�#�EP�M���
���E�P�MQ�M�#������I���_^[���   ;��������]�����������������������������������U����   SVW��@����0   �������EP�MQ�UR�EP����Q �BH�Ѓ�;��w���_^[���   ;��g�����]�������������������������������������U����   SVWQ��4����3   ������Y�M��} u�4�} t�EP�M�q���� �} t�EP�M�	����E�P�M�	��_^[���   ;��������]� �������������������������������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��B@��;��[���_^[���   ;��K�����]� ����������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M����   ��;������_^[���   ;��������]� ����������������������U����   SVWQ��4����3   ������Y�M���EP������   �M��BD��;��{���_^[���   ;��k�����]� ����������������������U����   SVWQ��4����3   ������Y�M�����P@��M��B`��;�����_^[���   ;�������]���������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P����Q@�B�Ѓ�;�����_^[���   ;�������]� �����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H@�Q�҃�;�����_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR����P@�M����   ��;�����_^[���   ;�������]� �������������������������������U����   SVWQ��4����3   ������Y�M���E P���E�$�MQ�UR�EP�MQ������   �M����   ��;������_^[���   ;��������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B@�HL�у�;��z���_^[���   ;��j�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M����   ��;������_^[���   ;��������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M��P\��;��z���_^[���   ;��j�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B@�M��Pp��;������_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP����Q@�M��Bh��;��~���_^[���   ;��n�����]� �������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ����B�M��Pp��;��
���_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M��B ��;�����_^[���   ;��t�����]� �������������������������������U����   SVWQ��(����6   ������Y�M���E�P����Q@�B�Ѓ�;������E�E�#Et�E��#E�E��	�E�E�E��E�P�M�Q����B@�H�у�;������_^[���   ;�������]� ��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR������   �M���D  ��;��A���_^[���   ;��1�����]� ����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B@�H�у�;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B@�H �у�;��J���_^[���   ;��:�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�����������������U����   SVW��@����0   �������j �EP����QD��Ѓ�;�����_^[���   ;��r�����]��������������������������������U����   SVW��@����0   �������j h�_ ����HD��҃�;�����_^[���   ;�������]��������������������������������U����   SVW��@����0   �������EPhO  ����QD��Ѓ�;�����_^[���   ;�������]�����������������������������U����   SVW��@����0   �������j �EP����QD��Ѓ�;��2���_^[���   ;��"�����]��������������������������������U����   SVW��@����0   �������j h:  ����HD��҃�;������_^[���   ;�������]��������������������������������U����   SVW��@����0   �������j h�  ����HD��҃�;��R���_^[���   ;��B�����]��������������������������������U����   SVW��@����0   �������EPh'  ����QD��Ѓ�;������_^[���   ;��������]�����������������������������U����   SVW��@����0   �������EP�MQ����BD��у�;��p���_^[���   ;��`�����]������������������������������U����   SVW��@����0   �������EPh2  ����QD��Ѓ�;������_^[���   ;��������]�����������������������������U����   SVW��@����0   �������j h�F ����HD��҃�;�����_^[���   ;�������]��������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��!����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��!����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��!����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��!����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;��!����E�     _^[���   ;�������]��������������������������������������U����   SVW��@����0   �������E�Q����B@�H�у�;������E�     _^[���   ;�������]��������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;��>���_^[���   ;��.�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;��^���_^[���   ;��N�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;������_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;��~���_^[���   ;��n�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;�����_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;��.���_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;��N���_^[���   ;��>�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;������_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;��n���_^[���   ;��^�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;������_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;�����_^[���   ;��~�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;��>���_^[���   ;��.�����]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B(�Ѓ�;������_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B�Ѓ�;��^���_^[���   ;��N�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H$�у�;������_^[���   ;��������]� �������������������������������������U���4  SVWQ�������M   ������Y�M���E�P������Q����BX�H�у�;��g����   ���}�E_^[��4  ;��H�����]� �����������������������������������U����   SVWQ��$����7   ������Y�M��M�������E�    �E�    �E�Pj�M��������u3���E�R��P�x��i���XZ_^[���   ;�������]Ð   ������   ��rp �������������������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����QD�B$�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ������;   ������Y�M���E�P�����Q����BX��у�;������U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;��p�����]� �������������������������������������������U����   SVWQ������;   ������Y�M���E�P�����Q����BX�H�у�;�������U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;�������]� ������������������������������������������U����   SVWQ������;   ������Y�M���E�P�����Q����BX�H�у�;��G����U��
�H�J�H�J�H�J�H�J�@�B�E_^[���   ;�������]� ������������������������������������������U����   SVWQ��$����7   ������Y�M��} u3��0�M�諢���E�    �E�E�E�Pj�M�貣����u3���   R��P�Ċ����XZ_^[���   ;��a�����]�    ̊����   ؊rp �����������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����HD�Q�҃�;������_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H �у�;��J���_^[���   ;��:�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H�у�;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H�у�;��J���_^[���   ;��:�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H�у�;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����BX�H�у�;��J���_^[���   ;��:�����]� �������������������������������������U����   SVW��@����0   �����󫡸��H\����;������_^[���   ;��������]��������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H0�у�;��j���_^[���   ;��Z�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�HH�у�;������_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H�у�;��j���_^[���   ;��Z�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�HD�у�;������_^[���   ;��������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q\�B�Ѓ�;��n���_^[���   ;��^�����]����������������������������U����   SVW��@����0   �������E�Q����B\�H�у�;������E�     _^[���   ;��������]��������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H\�Q8�҃�;��w���_^[���   ;��g�����]� ����������������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q\�B4�Ѓ�;������_^[���   ;��������]����������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q\�B�Ѓ�;�����_^[���   ;��~�����]����������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�EP�M�Q����B\�H`�у�;�����_^[���   ;��������]� �������������������������U����   SVWQ��4����3   ������Y�M���E�P����Q\�B�Ѓ�;�����_^[���   ;�������]����������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H@�у�;��*���_^[���   ;�������]� �������������������������������������U���  SVWQ�������B   ������Y�M��E�P�M�ߎ���}� |o�M������E�P�M�Ŏ���}� tU�E�    �	�E����E��E�;E�};�E�P�M虎���E�P�M荎���	�Eȃ��EȋE�;E��E�P�M�������봸   R��P� ������XZ_^[��  ;��%�����]�    �����   @�����   <�����   :�����   8�b a cnt level ��������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H�у�;��J���_^[���   ;��:�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H\�Q�҃�;������_^[���   ;�������]� ����������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H<�у�;��J���_^[���   ;��:�����]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�M�Q����B\�H �у�;������_^[���   ;�������]� �������������������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U�R����H\�Q$�҃�;��G���_^[���   ;��7�����]� ����������������������������������U����   SVWQ������?   ������Y�M�j �M裘���M��v����EȋE�P�M茘���E�    �	�E���E�E�;E�}3�E�P�M�Qh����U�R�M�趮���E�P�M�M����E�P�M�A����R��P�Ș����XZ_^[���   ;��]�����]�    И����   �����   �b a ��������������������������������������������������������������������U���,  SVWQ�������K   ������Y�M��}}�B  �E�E��E������E�E���EE�EȋE����EE�E��}�~�E���E�E�+E�E��1�EP�M�Q�U�R�M��j����E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��������}�Eԃ��EԋE��E���E�P�M�Q�U���M����;�������}�EP�M�Q�U�R�M�蕟�����U��������_^[��,  ;��o�����]� ����������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M������E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;��<�����}�Eԃ��EԋE��E���E�P�M�Q�U���M����;�������}�E�P�M�Q�U�R�M��7������U��������_^[��8  ;��������]� �����������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et.�E���E�M��U�E���E�M�U���E�M���_^[��]� ��������������������������������U���  SVWQ�������E   ������Y�M��} t�} t�} t�} u3��  kE E�E���E�P�MQ�U���M����;��V����Eȃ}� u
�E���   ��}� }3���   �E�   �E���E��E�;E���   �E�E����EԋE�E�E�E���E�P�MQ�U���M����;�������Eȃ}� uP�}� ~C�Eԃ��EԋE�E�E�E���E�P�MQ�U���M����;�������t�
��E��E�뷋E��#��}� }�Eԃ��E��	�Eԃ��E��G���3�_^[��  ;��[�����]� ������������������������������������������������������������������������������������������������������U���  SVWQ�������E   ������Y�M��} t�} t�} t�} u�E� ����3���  kE E�E���E�P�MQ�U���M����;��}����Eȃ}� u
�E��  ��}� }�E�     3��  �E�   �E���E��E�    �E�;E���   �E�E����EԋE�E�E�E���E�P�MQ�U���M����;�������Eȃ}� uS�}� ~C�Eԃ��EԋE�E�E�E���E�P�MQ�U���M����;�躾����t�
��E��E�뷋E���   ��}� }�Eԃ��E��	�Eԃ��E��D����}� ~�Eԃ��M���E�Mԉ�E�;M}F�E�M�M�M���E�P�MQ�U���M����;��0�����|h�a�8���9P�������E�8 ~I�E����MM�M���E�P�MQ�U���M����;��߽����h�a�8���?P�R�����3�_^[��  ;�賽����]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��u�EP�MQ�UR�M������Q�} uǅ0���   �
ǅ0���    ��0�����t�EP�MQ�UR�M��O�����EP�MQ�UR�M�赓��_^[���   ;��m�����]� ��������������������������������������������������������U���8  SVWQ�������N   ������Y�M��E���Eȃ}}�B  �E�E��E������E�E���EE�E��E����EE�E��}�~�E���E�E�+E�E��1�E�P�M�Q�U�R�M���|���E����E��}�u��   �E�+E�E��E�EԋEԃ��EE�E��E���;E���   �E����EԋE��E��Eԃ��EE�E��E�;E�}9�E�E�E���E�P�M�Q�U���M����;�������}�Eԃ��EԋE��E���E�P�M�Q�U���M����;��ݺ����}�E�P�M�Q�U�R�M���{�����U��������_^[��8  ;�觺����]� ������������������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E���E�M���M�U���U�E���Et4�E���E�Mf�f�U�E���E�M�Uf�f��Ef�M�f���_^[��]� ������������������������������������������U����   SVW��@����0   ������E;Et�&�} t �} t�} t�EP�MQ�UR������_^[���   ;��!�����]�������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��=����EP�M����.����EP�M���0�����EP�M���H�����E�_^[���   ;�萸����]� �������������������������������������������U���L  SVWQ�������S   ������Y�M��M��֎���M����ˎ���M���0������M���H赎�����x^�$���x^�$���x^�$�����������M����P�Q�P�Q�P�Q�P�Q�@�A���x^�$���x^�$����`�$������趫���M������P�Q�P�Q�P�Q�P�Q�@�A���x^�$����`�$���x^�$�������S����M���0���P�Q�P�Q�P�Q�P�Q�@�A����`�$���x^�$���x^�$����������M���H���P�Q�P�Q�P�Q�P�Q�@�A�E�_^[��L  ;��w�����]�������������������������������������������������������������������������������������������������������������������������������������U���  SVWQ�������C   ������Y�M��M��f����M����[�������b�$�����������E���������������P�� ����H������P������H������P����b�$�����迪���E���������������P�� ����H��$����P��(����H��,����P�E��@0    �E�_^[��  ;�������]�����������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��E� �E��E�@�E��E�@�E�_^[��]� ���������������������������U����   SVWQ��4����3   ������Y�M��E�_^[��]� �����������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�M�P;Quljj�M��͕����u��   �   k� �U���U���   �� �M���M�I��   ���M���M�I��   k� �U��B�   �}jj�M��a�����u�k�   k� �U���U���   �� �M���M�I��   ���M���M�I��   k��U���U�R��   k� �U��B�   �E�_^[���   ;�諲����]� ��������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �EP�M��I����E�_^[���   ;�������]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�_^[��]�����������������������������U����   SVWQ��4����3   ������Y�M��M�����_^[���   ;�������]������������������U����   SVWQ��4����3   ������Y�M��EP�M�� ����E�_^[���   ;�轰����]� ������������������������U���8  SVW�������N   ������j �M��՘���E�M�@8�YAX�U�E�JP�YH@�\��M�YA�U�E�JP�YH(�M�U�Q �YRX�\ʋE�YH0�X��M�U�I �YJ@�E�M�P8�YQ(�\ʋU�YJH�X��E��E�f.x^���Dz�M�?����E�  ��`�^E��E��E�M�@�YAX�U�E�JP�YH�\��M�YA0�U�E�J�YH8�M�U�Q�YR@�\ʋE�YHH�X��M�U�IP�YJ@�E�M�P8�YQX�\ʋU�Y
�X��YE��E��E�M�@�YA(�U�E�J �YH�\��M�YAH�U�E�J �YHX�M�U�QP�YR(�\ʋE�Y�X��M�U�IP�YJ�E�M�P�YQX�\ʋU�YJ�X��YE��E��E�M�@8�YA(�U�E�J �YH@�\��M�Y�U�E�J@�YH�M�U�Q8�YR�\ʋE�YH�X��M�U�I�YJ �E�M�P�YQ(�\ʋU�YJ0�X��YE��E��E�M�@8�YAX�U�E�JP�YH@�\��YE��E��E�M�@P�YA(�U�E�J �YHX�\��YE��E��E�M�@ �YA@�U�E�J8�YH(�\��YE��EċE�M�@@�YAH�U�E�JX�YH0�\��YE��E̋E�M�@X�YA�U�E�J(�YHH�\��YE��EԋE�M�@(�YA0�U�E�J@�YH�\��YE��E܋E�M�@0�YAP�U�E�JH�YH8�\��YE��E�E�M�@H�YA �U�E�J�YHP�\��YE��E�E�M�@�YA8�U�E�J0�YH �\��YE��E��   �u��}�ER��P� �����XZ_^[��8  ;��#�����]�   �����`   �mi ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��0����4   ������E�M� �Y�U�E�J�YH�X��M�U�I�YJ�X����$谖�����]��E�f.x^���Dz���x^�$�M������E�[��`�^E��E�E�@�YE���$�M�A�YE���$�U��YE���$�M�.����E_^[���   ;��ݩ����]���������������������������������������������������������������������������U����   SVW��@����0   ������E�@�YE���$�M�A�YE���$�U��YE���$�M�i����E_^[���   ;�������]��������������������������������������U����   SVW��@����0   ������E�M�@(�Y�U�XB�E�M�H@�YI�X��U�E�JX�YH�X����$�M�U�A �Y�E�X@�M�U�I8�YJ�X��E�M�HP�YI�X����$�U�E�B�Y �M�X�U�E�J0�YH�X��M�U�IH�YJ�X����$�M�3����E_^[���   ;�������]��������������������������������������������������������������������������������U����   SVW��@����0   ������E�M�@�\A���$�U�E�B�\@���$�M�U��\���$�M�a����E_^[���   ;�������]����������������������������������������������U����   SVW��@����0   ������E�M�@�XA���$�U�E�B�X@���$�M�U��X���$�M豚���E_^[���   ;��`�����]����������������������������������������������U����   SVW��@����0   ������E�M� �YA�U�E�J�Y�\����$�M�U�A�Y�E�M��YI�\����$�U�E�B�Y@�M�U�I�YJ�\����$�M�Ǚ���E_^[���   ;��v�����]����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E��M� �X�U���E��M�@�XA�U��B�E��M�@�XA�U��B�E�_^[��]� ��������������������������������������������U����   SVW��@����0   ��������E�$�?�����_^[���   ;��\�����]��������������������������U����   SVWQ��4����3   ������Y�M��E��x0 ��   �E��M� f/v�E��M�� �E��M�@f/Av�E��M�A�@�E��M�@f/Av�E��M�A�@�E�M�� f/Av�E��M��@�E�M��@f/A v�E��M�A�@ �E�M��@f/A(v�E��M�A�@(�`�E����M���Q�P�Q�P�Q�P�Q�P�I�H�U����E��
��J�H�J�H�J�H�J�H�R�P�E��@0   _^[��]� �����������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M������} ��   ��h0b�<���P�M��Q����B���   �у�;������U���E��8 u3��r�} tQ��h0b�<���
P�M��Q����B���   �у�;��ϡ���U��B�E��x u�E�P�0o����3���E��M�H�E��M�H�   �3�_^[���   ;�腡����]� ����������������������������������������������������������������U����   SVW��4����3   ������j�+  ���E��}� u3���E���H��;������_^[���   ;�������]�����������������������U����   SVWQ��(����6   ������Y�M�h�   �  ���E�}� t�E샸�    u3����EP�U�M����   ��;��k���_^[���   ;��[�����]� ��������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �  ���E�}� t�E샸�    u����/��EP�MQ�UR�EP�MQ�UR�E�M����   ��;�趟��_^[���   ;�覟����]� �������������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S  ���E�}� t�E샸�    u����/��EP�MQ�UR�EP�MQ�UR�E�M����   ��;������_^[���   ;�������]� �������������������������������������������������U���4  SVWQ�������  ������Y�M��x^�E��E�    j �M��ې��j �M��ѐ��j ��p����Đ���E��H�U�<�}���x  �} ��  ��P�����t��j ��0���茐���   k� �U��kM��U��A�E��Q�U��A�E��Q�U��A�EčE�P�   �� �U��kMQ������R�#p�������0����P��4����H��8����P��<����H��@����P��D����E�   �	�E܃��Eܸ   k� �U��B�U�;��   �E�P�M���E�k�MQ�����R�o������M��P�U��H�M��P�U��H�M��P�U��E�P��0���Q��(���R�������P��P����m����E���0����M���4����U���8����E���<����M���@����U���D����6������x^�$��H��������E��H������L����P��P����H��T����P��X����H��\����P��P���P��h���Q�n�����U��H��
�H�J�H�J�H�J�H�J�@�B����P����$�_����ݝ��������������X����$�������S_����ݝ����������f/������&  ����P����$�_����ݝ��������������`����$��������^����ݝ����������f/�������   �E��HP���x^�$����`�$���x^�$�������_���P������Q�������U����
�H�J�H�J�H�J�H�J�@�B�E��P�M��HQ������R�ʐ�����M��0���P�Q�P�Q�P�Q�P�Q�@�A��  ����X����$��]����ݝ��������������`����$��������]����ݝ����������f/�������   ����`�$���x^�$���x^�$�������@���P�E��HP�����Q�������U����
�H�J�H�J�H�J�H�J�@�B�E��P�M��HQ��(���R褏�����M��0���P�Q�P�Q�P�Q�P�Q�@�A�   ���x^�$���x^�$����`�$��H����|���P�E��HP��h���Q�%������U��0��
�H�J�H�J�H�J�H�J�@�B�E��HP�M��0Q������R��������M�����P�Q�P�Q�P�Q�P�Q�@�A�EP������Q�M������   ���}��E�    �	�E܃��E܋E�;E}�E��H�U܋E���E��ۋE���U�k�EP�MQ�����R���������M��P�U��H�M��P�U��H�M��P�UċE���U�kD�EP�MQ��0���R踕������M��P�U��H�M��P�U��H�M��P�U��E�    �	�E܃��E܋E��H�U�E�;���   �E܃��M��I�u��<�UЋE��k�UR�EP��P���Q�8��������p����H��t����P��x����H��|����P�U��@�E���p���P�M�Q�U�R�  ��ݝ�����������XE��E�E��E��M��M��U��U��E��E��M��M��U��Uċ�p����E���t����M���x����U���|����E��M��M��U��U�������E�R��P����e���XZ_^[��4  ;�訖����]� �I    ������   ������   ��p���   ��P���   ��0���   ��prev n v3 v2 v1 ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��8����2   ������E�M�@�\A�U�Y�E�M�H�\I�U�Y
�X��E�M�H�\I�U�Y
�X���8���݅8���_^[��]���������������������������������U����  SVWQ��<����q   ������Y�M��M��j���E�    �	�Ẽ��E̋E��M�;H�	  �E���U̍��p����u�ҋE���U̍��c����E�E��E��M��P;Qud�E�kMQ�U�kBEP��@���Q�Ee����P�U�kEP�M�kQUR��`���P� e����P������Q諈����P�M������c�E�kMQ�U�kBEP������Q��d����P�U�kBEP�M�kQUR������P�d����P������Q�F�����P�M�蹁��������E�P�MQ�ed�����ER��P� ��å��XZ_^[���  ;�������]� �   (�����   4�v ����������������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j �f   ���E�}� t	�E�x  u3����EP�U�M��B ��;��$���_^[���   ;�������]� �������������������������������U����   SVW��@����0   ������h���EPh_� �v����_^[���   ;�諐����]�������������������������U����   SVWQ��(����6   ������Y�M�j<�v������E�}� t	�E�x< u���EP�U�M��B<��;��6���_^[���   ;��&�����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�j8��������E�}� t	�E�x8 u3����E�M��P8��;�訏��_^[���   ;�蘏����]��������������������������������������U����   SVWQ��(����6   ������Y�M�jx�V������E�}� t	�E�xx u3����EP�MQ�U�M��Bx��;�����_^[���   ;�� �����]� �������������������������������������������U����   SVWQ��4����3   ������Y�M��M��jx���} �{  �} �q  ��h0b�D���P�M��Q����B���  �у�;��^����U���E��8 u3��0  �} ta�} t[��h0b�D���
P�M��Q����B���  �у�;������U��B�E��x u�M��w��3���   �E��M�H�Y�E��@   ��h0b�D���P�M��Q��R����H���  �҃�;�襍���M��A�E��x u�M��Tw��3��p�E��M�H�E��Q�U��B��P�M��R�EP��`�����} t&�E��HQ�U��B��P�M��QR�EP��`������   k� �U��B�U��   _^[���   ;��
�����]� ���������������������������������������������������������������������������������������������������������������������U����   SVWQ��4����3   ������Y�M��M��*v���} �.  �E�8 �"  �E�x �  ��h0b�@���P�M�Q��R����H���  �҃�;������M���E��8 u3���   �E�x tX�E�x tO��h0b�@���
P�M�Q��R����H���  �҃�;�賋���M��A�E��x u�M��bu��3��q�E��M�Q�P�E��M�Q�P�E��Q�U��B��P�M��R�E�Q��^�����E��x t'�E��HQ�U��B��P�M��QR�E�HQ��^�����   _^[���   ;�������]� ��������������������������������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�U�M��B��;��T���_^[���   ;��D�����]� �������������������������������U����   SVWQ��(����6   ������Y�M�jp�������E�}� t	�E�xp u3����EP�MQ�U�M��Bp��;������_^[���   ;�谉����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jT�f������E�}� t	�E�xT u���E�M��PT��;��*���_^[���   ;�������]����������������������������������������U����   SVWQ��4����3   ������Y�M��E����   @t�����E�� %���3ҹ   ���_^[��]��������������������������������U����   SVWQ��(����6   ������Y�M�j4�f������E�}� t	�E�x4 u������EP�MQ�U�M��B4��;�����_^[���   ;�������]� ������������������������������������������U����   SVWQ��(����6   ������Y�M��} |�E��8 u����<�E�    �	�E���E�E��M�;H}�E���U���uW��;Eu�E���Ѓ��_^[���   ;��]�����]� ����������������������������������������U����   SVWQ��4����3   ������Y�M��E�P�|T�����E���P�mT�����E��@    �E��@    _^[���   ;��͆����]���������������������������U����   SVW��(����6   ������E�8 u�>j�������E��}� u�)�E��M��E�P�M��Q�҃�;��R����E�     R��P�������XZ_^[���   ;��(�����]Ð   �����   �i ����������������������������������������������U����   SVWQ��(����6   ������Y�M�j\��������E�}� t	�E�x\ u���E�M��P\��;�芅��_^[���   ;��z�����]����������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �3������E�}� t�E샸�    u���EP�U�M����   ��;�����_^[���   ;��݄����]� ����������������������������������������U����   SVWQ��(����6   ������Y�M�jh�������E�}� t	�E�xh u�(��EP�MQ�UR�EP�MQ�U�M��Bh��;��F���_^[���   ;��6�����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�j(��������E�}� t	�E�x( u3����E�M��P(��;�踃��_^[���   ;�訃����]��������������������������������������U����   SVWQ��(����6   ������Y�M�jP�f������E�}� t	�E�xP u3����E�M��PP��;��(���_^[���   ;�������]��������������������������������������U����   SVWQ��$����7   ������Y�M��M��R����E�E�M���R����$�����$�������$�����$���w}��$����$� ��E� ����E� ����\�E�M���E�M�Q��E�E�M�Q��E�M�Q��-�E�M�Q��E�M�Q���E�M�Q��E�M��_^[���   ;�������]� �I ��������������������������������������������������������������������������������������U����   SVWQ������9   ������Y�M��E� �E�    �	�E����E��E��M�;H}3�E���U����DQ��;Eu�]�E���U����Z�����؈]���E���_^[���   ;�������]� ���������������������������������������������U����   SVWQ��(����6   ������Y�M�j$��������E�}� t	�E�x$ u2����EP�U�M��B$��;�脀��_^[���   ;��t�����]� �������������������������������U����   SVWQ��(����6   ������Y�M�jL�6������E�}� t	�E�xL u3����E�M��PL��;�����_^[���   ;�������]��������������������������������������U���L  SVWQ�������S   ������Y�M��E��x0 ��   ����^�$�E���P�M�Q������R�n�����P������P�Ϗ�����M���P�Q�P�Q�P�Q�P�Q�@�A�EP�M���Q������R�yQ�����M���P�Q�P�Q�P�Q�P�Q�@�A�{���x^�$������Ht���E������������P�� ����H��$����P��(����H��,����P�E�M���P�Q�P�Q�P�Q�P�Q�@�A_^[��L  ;��d~����]� �����������������������������������������������������������������������������������������������U���$  SVWQ�������I   ������Y�M��M���Y���E�    �	�E����E��E��M�;H��   �E���U�����Z����u�ҋE���U����M����E�E��E�kMQ�M��\���E�kHMQ�M��\���E�kHMQ�M��\���E��M��P;Qt�E�kHMQ�M��t\���[����EP�MQ�M���?��R��P�0�貐��XZ_^[��$  ;���|����]�    8�����8   D�mm �������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j,�v������E�}� t	�E�x, u3����E�M��P,��;��8|��_^[���   ;��(|����]��������������������������������������U����   SVWQ������9   ������Y�M��E�    �E�    �	�E����E��E��M�;H} �E���U�����K�����t	�E���E��̋E�_^[���   ;��{����]�����������������������������������U����   SVWQ������9   ������Y�M��E�    �E�    �	�E����E��E��M�;H}�E���U����bX����t	�E���E��͋E�_^[���   ;���z����]������������������������������������U����   SVWQ������9   ������Y�M��E�    �E��x|�E��8 u3��?�E�    �	�E����E��E��M�;H}�E���U����H����t	�E���E��͋E�_^[���   ;��1z����]�����������������������������������������������U����   SVWQ��(����6   ������Y�M��E�E��	�E���E�E��M�;H}!�E���U����G����t�E�+E����˃��_^[���   ;��y����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�jX�F������E�}� t	�E�xX u���E�M��PX��;��
y��_^[���   ;���x����]����������������������������������������U����   SVWQ��4����3   ������Y�M��E�� %    _^[��]�����������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3����EP�MQ�U�M����   ��;��x��_^[���   ;��x����]� ����������������������������������U����   SVWQ��(����6   ������Y�M�j��������E�}� t	�E�x u3�� ��EP�MQ�UR�E�M��P��;��|w��_^[���   ;��lw����]� ���������������������������������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    _^[��]��������������������������������U����   SVWQ��(����6   ������Y�M�jl�������E�}� t	�E�xl u3�� ��EP�MQ�UR�E�M��Pl��;��lv��_^[���   ;��\v����]� ���������������������������������������U����   SVWQ��(����6   ������Y�M�jt�������E�}� t	�E�xt u3����EP�MQ�U�M��Bt��;���u��_^[���   ;���u����]� �������������������������������������������U����   SVWQ������9   ������Y�M��M��]E���E�M��E���E��E;E�t	�}���u�E;E�t	�}���u�^�}���t�E�E��}���t�E�E�}��t�E�M����E����   �ыE����E���   @�M����   �M��_^[���   ;���t����]� ���������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j`�f������E�}� t	�E�x` u3����EP�MQ�U�M��B`��;�� t��_^[���   ;��t����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�jD��������E�}� t	�E�xD u3����EP�U�M��BD��;��s��_^[���   ;��ts����]� �������������������������������U����   SVWQ��(����6   ������Y�M�j0�6������E�}� t	�E�x0 u3����EP�U�M��B0��;���r��_^[���   ;���r����]� �������������������������������U����   SVWQ��(����6   ������Y�M�jH�������E�}� t	�E�xH u���EP�U�M��BH��;��fr��_^[���   ;��Vr����]� ���������������������������������U����   SVWQ��(����6   ������Y�M�h�   �������E�}� t�E샸�    u3��#��EP�MQ�UR�E�M����   ��;���q��_^[���   ;��q����]� ����������������������������������������������U����   SVWQ��(����6   ������Y�M�h�   �c������E�}� t�E샸�    u3����EP�MQ�U�M����   ��;��q��_^[���   ;��q����]� ����������������������������������U����   SVW��@����0   ��������E�$��+ ��_^[���   ;��p����]��������������������������U����   SVWQ��(����6   ������Y�M��M��@���E�}��u3��
�   �M���_^[���   ;��-p����]���������������������������U����   SVWQ��(����6   ������Y�M�jd��������E�}� t	�E�xd u3����EP�MQ�U�M��Bd��;��o��_^[���   ;��o����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M�j�V������E�}� t	�E�x u3����EP�U�M��B��;��o��_^[���   ;��o����]� �������������������������������U����   SVWQ��(����6   ������Y�M�j@��������E�}� t	�E�x@ u���EP�U�M��B@��;��n��_^[���   ;��vn����]� ���������������������������������U����   SVWQ������<   ������Y�M��E�    �	�E���E�E��M�;H}�E���U��%����M���M�����E�    �	�E���E�E��M�;H}{�E���U��%   �ud�E���U���=���EԋE���E��	�E����E��E��M�;H}2�E���U����z=��;E�u�E���U���   ��M���M�����q���_^[���   ;��Jm����]������������������������������������������������������������������������U����   SVWQ��(����6   ������Y�M�j|��������E�}� t	�E�x| u3����EP�U�M��B|��;��l��_^[���   ;��l����]� �������������������������������U����   SVWQ��(����6   ������Y�M�h�   �S������E�}� t�E샸�    u3��'��EP�MQ�UR�EP�U�M����   ��;���k��_^[���   ;���k����]� ������������������������������������������U����   SVWQ��(����6   ������Y�M�j�������E�}� t	�E�x u3����EP�U�M��B��;��dk��_^[���   ;��Tk����]� �������������������������������U����   SVW��(����6   ������} t�E�8 t�E� �Pj�EP�A�����E��}� u3��5�M���2���E�}� u3�� �} t�E�M��E�M;H~3���E�_^[���   ;��j����]������������������������������������������U����   SVW��@����0   ������E�M��E�M�H�EPj�MQ�r����_^[���   ;��j����]����������������������������U����   SVW��@����0   ������   _^[��]�����������������������U����   SVW��4����3   ������E��M��E�M���E�M��_^[��]������������������U����   SVWQ��4����3   ������Y�M��M���S���E�� $c�E��M�H�E�_^[���   ;��i����]� ��������������������������U����   SVWQ��4����3   ������Y�M��E�� �b�M�����p���M�����p���E��@    �M��7Z���E�_^[���   ;��h����]��������������������������������������U����   SVWQ��4����3   ������Y�M��E�� �b�E��@    �E��@    �E�_^[��]�����������������������U����   SVWQ��4����3   ������Y�M��E�� �b�M���(��_^[���   ;���g����]�������������������������U����   SVWQ��4����3   ������Y�M��E�� �b�M��m���M����s���M����ws��_^[���   ;��Ug����]�����������������������������������U����   SVWQ��4����3   ������Y�M��E�� �b�M���@��_^[���   ;���f����]�������������������������U����   SVWQ��4����3   ������Y�M��M���5���E��t�E�P�az�����E�_^[���   ;��}f����]� ������������������������U����   SVWQ��4����3   ������Y�M��M��Q���E��t�E�P��y�����E�_^[���   ;��f����]� ������������������������U����   SVWQ��4����3   ������Y�M��M���q���E��t�E�P�y�����E�_^[���   ;��e����]� ������������������������U����   SVWQ��4����3   ������Y�M��E��M��P;Qu�M��:]����u3��&�E��H�U��B�U���E��H���U��J�   _^[���   ;��e����]� �����������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E����M�A�E�M��Q�P�E��H�U�Q�E��M�H_^[��]� ���������������������������������U����   SVWQ��4����3   ������Y�M��E��@    �E����M��A�E����M��A�E��@    _^[��]���������������������������U����   SVWQ��4����3   ������Y�M���EP�MQ�U��B�Ѓ�;��c��_^[���   ;��c����]� ���������������������������U����   SVWQ��(����6   ������Y�M��M�C$���E�M��Q�P�E�M��Q�P�E�    �	�E���E�E��M�;H}�E��H�U��P�M��w����u3���͸   _^[���   ;���b����]� ��������������������������������������U����   SVWQ������9   ������Y�M��E��x u�E��H�M��%�E��x t�E��H�U�J�M���E��H��M��}� u3��]��h�b�H���P�M���Q�U��BP����Q��  �Ѓ�;�� b���E�}� u3���E��M�H�E��M��H�   _^[���   ;���a����]����������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�    �	�E���E�E��M�;H}�E��H�U��;Eu�E���ԃ��_^[��]� ����������������������������U���   SVWQ�� ����@   ������Y�M��M��h���E��}� tm�M��A���E�}� tM�E��������������������� t%��j��������������;��`���� ����
ǅ ���    �E�    �E�E�덋M��R��_^[��   ;��v`����]����������������������������������������������������U����   SVWQ��4����3   ������Y�M��E���P�-�����E��@    �E��@    �M��A    _^[���   ;���_����]�����������������������������U����   SVWQ������9   ������Y�M��E�    �M��?g���E���M��'@���E��}� t�E���E���E�_^[���   ;��Y_����]���������������������������������������U����   SVWQ��0����4   ������Y�M��E����M�9At�U��B��0����
ǅ0���    ��0���_^[��]���������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H}�E��H�U���3�_^[��]� �������������������U����   SVWQ������<   ������Y�M��E�    �M���e���E��}� tZ�E쉅����M������U���U싅���;����uǅ���   �
ǅ���    ����� t�E���M��v>���E��3�_^[���   ;��]����]� ���������������������������������������������������U����   SVWQ��0����4   ������Y�M��E��x t�M��Q�z t�E��H��0����
ǅ0���    ��0���_^[��]������������������������������������U����   SVWQ��(����6   ������Y�M��E��M;H~	�E��H�M�} }�E    �E��M��P;Qu�M��T����u3��Z�E��H�M��	�E���E�E�;E~�E��H�U��B�U�u�L�����ԋE��H�U�E���E��H���U��J�   _^[���   ;��3\����]� ��������������������������������������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E�M��Q�P�E����M�A�E��H�U�Q�E��M�H_^[��]� ���������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E��M�Q�P�E�M��H�E��M�H�E��H�U��Q_^[��]� ������������������������������������U����   SVWQ��(����6   ������Y�M��E�E�E��M�Q�P�E�M��H�E��M�H�E��H�U��Q_^[��]� ������������������������������������U����   SVWQ��(����6   ������Y�M��E;E}	�E���E�} |$�E��M;H}�} |�E��M;H}�E;Eu�/�E��H�U���E�EP�M���m����t�EP�M�Q�M��HB��_^[���   ;���Y����]� �������������������������������������������U����   SVWQ��(����6   ������Y�M��E��H��Q�M��R?���E�}� t�E��H��Q�M��"m���E�_^[���   ;��<Y����]��������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|3��E�E��H���U��J�	�E���E�E��M;H}�E��H�U��B�U�u�L����Ѹ   _^[��]� ������������������������������������������U����   SVWQ��4����3   ������Y�M��EP�M��[��P�M��
l��_^[���   ;��'X����]� ����������������������������������U����   SVWQ��4����3   ������Y�M��E��x t;�E��x t2�E��H�U��B�A�E��H�U��B�A�E��@    �M��A    _^[��]�����������������������������������U����   SVWQ������9   ������Y�M��M���^���E��}� t�M���7���E�M���0���E�E���_^[���   ;��W����]������������������������������U����   SVWQ��4����3   ������Y�M��E��@    _^[��]�����������������������������U����   SVWQ��$����7   ������Y�M��EP�M��F:��j�E��HQ�U��BP�MQ�M��	`��R��P��	��i��XZ_^[���   ;��3V����]� ��   �	����   
sort �����������������������������������U����   SVWQ��4����3   ������Y�M��} |�E��M;H|3���E��H�U�E���   _^[��]� ���������������������������U����   SVWQ��4����3   ������Y�M��E��M;H}�EP�MQ�M��R���#�E��H;M}j �M��j����EP�M���i��_^[���   ;��U����]� ���������������������������������������U����   SVWQ��$����7   ������Y�M��EP�M��8��j�E��HQ�U��BP�M�����R��P���4h��XZ_^[���   ;��wT����]� ��   �����   �sort ���������������������������������������U����   SVWQ��4����3   ������Y�M��} |$�E��M;H}�} |�E��M;H}�E;Eu�"�E��H�U��P�M��Q�E��Q������_^[���   ;��S����]� �����������������������������������������U����   SVW��@����0   ������h���EPh�f �9����_^[���   ;��;S����]�������������������������U����   SVW��4����3   ������j�{������E��}� t	�E��x u3����EP�MQ�U��B�Ѓ�;���R��_^[���   ;��R����]�����������������������������������U����   SVW��4����3   ������j��������E��}� t	�E��x u����0��E P�MQ�UR�EP�MQ�UR�EP�M��Q�҃�;�� R��_^[���   ;��R����]����������������������������������������������U����   SVW������<   ������j�;������E��}� t	�E��x uǅ��������M����������E�E8P�M4Q�U0R�E,P�M(Q���̍UR��Z���EP�M��Q�҃�4�� ����M����� ���_^[���   ;��6Q����]����������������������������������������������������U����   SVW��4����3   ������j�[������E��}� t	�E��x u3����EP�M��Q�҃�;��P��_^[���   ;��P����]���������������������������������������U����M��L��   ��Au,�E�    �	�U����U��}�}kE���P�vX�����݋E���]��������������������U��Q�M��E��M��U��: uj�S������E��8}�M�k����R��X�����E���]� �����������������������U��Q�M��E��     �M��9 uj��������   k� ��P�~X�����E���]��������������������������������U����M��L������Iy,�E�    �	�U����U��}�}kE���P��B�����݋�]�������������������������U��Q�M��E��8 uj�M������M��9}�U�k��P��<������]����������������������U��Q�L��   ��Au,�E�    �	�U����U��}�}kE���P�V�����݋�]����������������������������U��Q�L������Iy,�E�    �	�U����U��}�}kE���P��A�����݋�]������������������������������U��   k� ����Q��V����]���������������������U��} uj�������E���M��Uk��P�V����]���������������������������U��} uj�������E��k�����Q�;V����]������������������U��Ek����Q�N;����]�������U��} uj�K������E��k�����Q�;����]������������������U���%��]�������U��EP�MQ�UR��#����]��������U��EPh�Yj �MQ�URj��������u�]�������������������������U��} u�EP�MQhH]�v#����]�����������������U��Q�M��E���]�������������������U��Q�M��EP�M��T���M��dh�E���]� �����������U����M��E�phj�E�P�M��T���M��dh�E���]�������������������U��Q�M��EP�M��2T���M���h�E���]� �����������U��Q�M��M��>���E�� �h�E���]� ���������������U��Q�M��EP�M��w;���M���h�E���]� �����������U��Q�M��EP�M���B���M���h�E���]� �����������U��Q�M��EP�M��;���M���h�E���]� �����������U��Q�M��EP�M��{B���M���h�E���]� �����������U��Q�M��EP�M��S���M���h�E���]� �����������U��Q�M��EP�M���"���M���h�E���]� �����������U��Q�M��EP�M��W:���M���h�E���]� �����������U��Q�M��EP�M��A���M���h�E���]� �����������U��Q�M��EP�M��/���M���h�E���]� �����������U��Q�M��EP�M��5���M���h�E���]� �����������U��Q�M��EP�M��V/���M�� i�U��E�H�J�E���]� ���������������U��Q�M��EP�G[����P�M�����M�� i�U��E�B�E���]� �������������������������U��Q�M��E�� dh�M��Y(����]���������������������U��Q�M��M��2(����]��������������U��Q�M��M��A+����]��������������U��Q�M��M��!+����]��������������U��Q�M��M���'����]��������������U��Q�M��M���*����]��������������U��Q�M��M��1����]��������������U��Q�M��M������]��������������U��]������������U��Q�M��M�����E��t�M�Q�M[�����E���]� ��������������������U��Q�M��M��{N���E��t�M�Q�[�����E���]� ��������������������U��Q�M��M��\U���E��t�M�Q��Z�����E���]� ��������������������U��Q�M��M������E��t�M�Q�Z�����E���]� ��������������������U��Q�M��M��q)���E��t�M�Q�MZ�����E���]� ��������������������U��Q�M��M��+9���E��t�M�Q�Z�����E���]� ��������������������U��Q�M��M���$���E��t�M�Q��Y�����E���]� ��������������������U��Q�M��M���E���E��t�M�Q�Y�����E���]� ��������������������U��Q�E�E��}�ws�M��$��i�g��i�`��i�Y�hj�R��j�K� k�D�xk�=��k�6�@l�/��l�(�Pm�!��m��Xn��o��(o��Ho��]Ú����������������������������������������������������������������������U����M��P��h�=�E�P�=����]�����������������U���j �M�����h?�E�P��<����]���������������U����EP�M��0
��h�=�M�Q�<����]�������������U����EP�M��-��h8>�M�Q�o<����]�������������U����EP�M��G=��h�>�M�Q�?<����]�������������U����EP�M���L��h�>�M�Q�<����]�������������U����EP�M���=��hT?�M�Q��;����]�������������U����EP�M����hT<�M�Q�;����]�������������U��Q�M���h��]�����������������U����".���E�h�   h�ojjh   � �����E�}� t h   ���P�E�P�m�����E�   �����E��E�    ����   �� ��U��}� t�E�P�6�����E��M�U���E�A�U��Q�E��A�E��]�������������������������������������������������������U���$�} u����   ���U��*-���E���E�H�M��U��E܃}� u�}A|�}Z	�M�� �M�E�  �}   s:�} u�UR�E9������u�E�i  ��E�H�U�Q��u�E�M  �} u"�����M�����   ���P% �  �E��4�M�����   �U�B�H�� �  t	�E�   ��E�    �U�U�}� tN�E��%�   �   k� �D��   �� �M�L��   ��U�}�s��#E���E��D� �E�   �2�   k� �E�D��E�   �}�s���D���M��D� �E�   j�U�Rj�E�P�M�Q�U�Rh   �E�Pj ��>����$�E�}� u�E�6�}�u�   k� �D��!��   �� �D��   k� �L������]���������������������������������������������������������������������������������������������������������������������������������U���$�} u����   ���U��*���E���E�H�M��U��E܃}� u�}a|�}z	�M�� �M�E�  �}   s:�} u�UR��=������u�E�i  ��E�H�U�Q��u�E�M  �} u"�^���M�����   ���P% �  �E��4�M�����   �U�B�H�� �  t	�E�   ��E�    �U�U�}� tN�E��%�   �   k� �D��   �� �M�L��   ��U�}�s��B���E��D� �E�   �2�   k� �E�D��E�   �}�s��B���M��D� �E�   j�U�Rj�E�P�M�Q�U�Rh   �E�Pj �k<����$�E�}� u�E�6�}�u�   k� �D��!��   �� �D��   k� �L������]���������������������������������������������������������������������������������������������������������������������������������U��} tj �M�%���EP�G����]����������������U��Q�M��E��     �M��A �UR�M������E���]� ��������������������U��Q�M��E��M��U��E�B�E���]� ���������������U��j�h��d�    PQ���3�P�E�d�    �M�j�M������E�    �E�� $p�M��A    �U��E�H�J�U��E�H�J�U��E�H�J�M���1��P�M�������E��UR�E�P�P'�����E������E��M�d�    Y��]� ������������������������������������������������������������U��j�h(�d�    PQ���3�P�E�d�    �M�j�M������E�    �E�� $p�M��A    �U��B    �E��@    �M��U�Qh4p�M����2
���E������E��M�d�    Y��]� ����������������������������������������������U��Q�M��E��M��E���]� ��������U��Q�M��E���]� ����������������U��Q�M��E��H�U���J�P��P��������]����������U����M��=x� t!�x��E��M���x��E�P�������֋�]��������������������������U��Q�M��E�� $p�M�Q��)�����M�����;���M�������]��������������U��EP�����]����������������U����M��E��;Mtv�M�����} th�U�U��E����t�U����U���E����E��M�+M�M�h-  h<pj�U�R��������M���U��: t�E�P�MQ�U��P�������E���]� ����������������������������������������������U��Q�M��M���'���E��t�M�Q�L�����E���]� ��������������������U��Q�M��M��E���E��t�M�Q�q�����E���]� ��������������������U����M��E��8 t
�M���U��	�E����E��E���]����������������������U����M��E��8 u	�E�   ��E�    �E���]�������������������������U��j�hh�d�    P�����3�P�E�d�    �1���E�j8h�o�E�Pj��K�����E��E�    �}� t�MQ�x�R�M��2���E���E�    �E�E��E������M�x��M�d�    Y��]�������������������������������������������U�졄�]�������U��j�h��d�    P�����3�P�E�d�    �E�    j �M������E�    �o=���E��}� ��   j ������E��E�P�8�����M��A?   h8p�M�������U������������B��h��j�������E��E��}� t���Q�M��;E���E���E�    �U�U��E� �E��t�M���M��B���E������M��J3���E��M�d�    Y��]�����������������������������������������������������������������������������U��j�h��d�    P�����3�P�E�d�    j �M��k���E�    �E�H�M��}� vB�U����U��E�H�U��<� t(�E�H�U����M�Q�M�� ���P��P�����븋E�HQ��?�����E������M��G2���M�d�    Y��]�������������������������������������������������������������U���j j �Z3�����E��}� u	�E��Q��E��E��M�Q�M��$����} t�URj �3�����E�} u	�E�4p��E�E�M�Q�M��,�c����]�����������������������������������������U��M��$�2������u�M��$���Pj �2����]��������������������U��j�h+�d�    P�����3�P�E�d�    �-���E�h�   h�o�E�Pj �	�����E��E�    �}� t�MQ�M���6���E���E�    �U�U��E������E�M�d�    Y��]�������������������������������������U��j�h{�d�    P�����3�P�E�d�    ��,���E�h�   h�o�E�Pj �\�����E��E�    �}� t�MQ�M��]���E���E�    �U�U��E������E�M�d�    Y��]������������������������������������U�������u���h`.�)�����M���]��������������������U��j �#�������]�������������U��Q�E�    j �#����j������P�M��@���E����E��E��]�������������������������U��Q�E��M��}� t�U���M��P��P�6������]���������������������U��Qj �M��l��h�����������    �M��.����]����������������U��Q�EP�MQ�U�P�MQ��������E��}� u�U���E���]��������������U��E�Q�UR�;����]����������U��EP�MQ�UR�EP�E����]��������������������U��EP�MQ�UR�EP�D����]��������������������U��pp]�������U��Q�   k� ���r�M��	�U����U��E��x t�M��;Uu�E��@���3���]������������������������������U��Q�   k� ��xp�M��	�U����U��E��x t�M��;Uu�E��@���3���]������������������������������U��} t�EP�n:����]����������U��} t�EP�N:����]����������U���j�M��Z���E�@    �M�Q���U��E�M��H�}�s&�U�B�<��� t�M�Q����;Eu�뿋M�Q�E�����M�Q�����M�Q�����M��/,����]������������������������������������������������U����M��E��H,�M���U���E��}� t�M��QR�E�P�MQ�U��B�Ѓ��֋�]� ����������������������������U��Q�E�x v*�M�Q����,�E��M�Q�E������M���~��M�����U�B0P��������]�������������������������������U����M�j �M��: ���E��H(�M���U��U��}� t�E���M��U�R� �����ދE��@(    �M��Q,�U���E�E�}� t�M��U�E�P�8�����ދM��A,    ��]��������������������������������������������U����E�    �E���E��M��   �M�U��@t	�E���E�M��t	�U���U�E%;����E�E�    �	�M����M��U��<�h� t�E���h�;Mt�ًU��<�h� u	3��   �x�}� t5�E��
t-�MQj �UR�������E��}� t�E�P�^����3��l�=�}� t�M�Q�F������t3��P�!�UR�E�P�MQ������E��}� u3��-�}� tjj �U�R��������u�E���E�P������3���]�����������������������������������������������������������������������������������U����E�    �E���E��M��   �M�U��@t	�E���E�M��t	�U���U�E%;����E�E�    �	�M����M��U��<��� t�E�����;Mt�ًU��<��� u	3��   �x�}� t5�E��
t-�MQj �UR�;������E��}� t�E�P������3��l�=�}� t�M�Q�������t3��P�!�UR�E�P�MQ��������E��}� u3��-�}� tjj �U�R��������u�E���E�P�`����3���]�����������������������������������������������������������������������������������U��EP�MQ�UR�Y�����]��������U��EP�MQ�UR�v.����]��������U��EP�MQ�UR������]��������U��EP�M��P�R�EP������]�����������������U��EP�M��ĀR�EP�)����]�����������������U��EP� ]������������������U��j h�  �EP�Y����]���������U��EP�  ]������������������U��EP� ]������������������U��Q�E�8u�F�   �U�
�M��}� u�U�E�    �%�}�u�M�   ��U�:tj�@&�������]�������������������������U����M�=X�
s6�X������M��X����X��E�P� �E��}� t�U�����]���������������������U��=X� u�����$�X����X��MQ� �X�����]������������������������U��]����������U��EP�M�.��]����������������U��Q�EP�M���
��P�MQ�M���
��P�	8������]�����������������������U��Q�EP�MQ��7�����Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ������Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ������Ѕ�u	�E�   ��E�    �E���]���������������U��} t�EP�>1����]����������U��} u�EP�MQhH]�������]�����������������U��]������������U��E;EtE�MQ�UR�EP�������MQ�UR�EP�������M;Ms�UR�EPh�]�T�����]�������������������������������U��Q�EP�MQ�J�����E��U��U���]����������������U��Q�EP�M�Q���������P�MQ�UR�EP�MQ�������]���������������������������U��Q�EP������E��M�Q�UR�EP�MQ�UR�EP�MQ��������]���������������������U��Q�E�E��	�M����M��U����t�M���E;�t�݋E�+E��]������������������������U��j�h��d�    P��D���3ŉE�VP�E�d�    �E�    �	�E����E��MM����t'�EE���   k� �U�;�u	�M���M��j �UR�M��R����E�    �E������E�   ��Eă��EċM�����E������E� �E�    �E�    �	�Mȃ��MȋU�;U�#  �	�EЃ��EЋMM����t�EE���   k� �U�;�t�̋M�Q�M���������t�E�P�M������MЉM��   �U�UĉUЋEE���   k� �U�;�t�MM����u.�}�s�EĉE���E�   �M�Q�M��Y����U���EȉE��[�MQ�UR���������u�MM��1�M������;�t(�}�s�EĉE���E�   �M�Q�M�������U����E�������Eυ�t�MQ�UR�.��������t��v����M��M��E������M��
����E��M�d�    Y^�M�3������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M��EPj �   k� �E��R�������M��A�URj �   k� �U�B�Q�Y������U��B��]�4 ����������������������U��Q�E���]������U��E]���������U����EP���������E�h�  h�����P�M�Q�������E��U��U�E�E���M����M��U����U��E���E�}� v�M��U���ӋE��]����������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��;����E�    �d��E�\��X����E�M�Q�M����E�}� t�n�}� t�U��U��`�EP�M�Q����������uh|]�M��K���hH=�U�R����.�E��E�M��d��U��U�E��M�B�ЋM�Q�#�����U�U��E������M������E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h(�d�    P��$���3�P�E�d�    j �M�������E�    �h��E�`������E�M�Q�M�i���E�}� t�n�}� t�U��U��`�EP�M�Q�~�������uh|]�M�����hH=�U�R�O���.�E��E�M��h��U��U�E��M�B�ЋM�Q��!�����U�U��E������M�����E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hX�d�    P��$���3�P�E�d�    j �M������E�    �l��E���������E�M�Q�M�)���E�}� t�n�}� t�U��U��`�EP�M�Q��������uh|]�M������hH=�U�R����.�E��E�M��l��U��U�E��M�B�ЋM�Q� �����U�U��E������M��W���E܋M�d�    Y��]��������������������������������������������������������������������������U��Q�M��E��     3ɋU�f�J�E���]�����������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M�������E�    �M�� ��UR�M�������E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��l����E�    �M��H��UR�M�����E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M�������E�    �M�����UR�EP�M��>����E������E��M�d�    Y��]� ����������������������������������U��Q�M��M�������]��������������U��Q�M��E��  ��M��������]���������������������U��Q�M��E�� H��M�������]���������������������U��Q�M��E�� ���M�����M��j�����]�������������U����M��E�;EtZ�M�Q�M���P�U�R�M����P�z���������t%3�t!j j�M�������U�R�M�s��P�M��J���EP�M�������E���]� ��������������������������������������������U����M��E��x t2�MQ�U��J�H
���E��C���E�E�P�M�Q�y�����Ѕ�t�E�� �E���]� �����������������������������U��Q�M��E��H;Msh�  hXohd��k������M��� ��E��]� ����������������������U��Q�M��E��H;Msh�  hXohd��������M��X��E��]� ����������������������U��Q�M��E��H��u�M�������U��: uh�  hЄh8��������E��@��]������������������������������U��Q�M��E���]�������������������U��Q�M��E��8 uh  hЄh���N������M�����E���]����������������������������U��Q�M��E���]�������������������U��Q�M��EP�M��>�����]� �������U��Q�M��EPj�M��������]� ��������������������U��Q�M��M��;����E��t�M�Q�������E���]� ��������������������U��Q�M��M��x����E��t�M�Q��������E���]� ��������������������U��Q�M��M������E��t�M�Q�������E���]� ��������������������U��Q�M��EP�MQ�U�R�F�������]� ���������������U��Q�M���]� ���U����E�E�M��%�U���U�E�� t�M��+�U���U�E��t�M��#�U���U�E�� .�M���M�U��*�E���E��M��t�U�E��M���M�U�� 0  �U��E��tP�}�    u�E�f�.�}� 0  u�E�A��}�   u�E�E��E�G�M��M��U��U��E�M���U���U��N�}�    u�E�f�.�}� 0  u�E�a��}�   u�E�e��E�g�E��E��M��M��U�E���M���M�U�� �E��]����������������������������������������������������������������������������������U��j�h6�d�    P���   ���3ŉE�SP�E�d�    h`  h���EP������}0 v�M ���+t�E ���-u	�E�   ��E�    �U��U��M����% 0  = 0  tǅ|���X��Jǅ|���\��E���;E0w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M���|���R�   k� M Q�"!�����E�f�`�f�U��6����   k� � �   k� ��T��   k� �T�R�   k� M Q�� �����E���`���R�M������l�����l�����\����E�    ��\���Q��������E��E�������`����=���j0�M�� ���E�j �U0R�M��/����E�   j �M��3���P�E E0P�   k� U R�M��'�����p���P�M�������d�����d�����h����E���h���R�"�����E��E���p��������E�P�M������E��M��M
���E��M$�M��U�;U0u �E�E��E��M�Q�U$R�E�P�M��"���c�M�M��M��U�R�E,P�M�Q�M���!���U�R�E(P�M���Q�M���!���M��K����؋U�R�M��<�����E�P�M$Q�U�R�M��!��j �M��~����E��E����tY�U����~O�M���E�+E�;�s?�M���E�+E��M�Qj�U�R�M��S!���   �� �M����~	�E����E�뜍M�������E0�M�V����t�����x�����x��� |(	��t��� v�M�.��;E0v�M�!��+E0�E���E�    �M��M��M���%�  �E��}�@ty�}�   tp�U�R�EP�MQ�UR��<���P�MQ�"�������@�U�E�E�    �M�Qj �M������P�UR�EP��T���Q�UR��������P�M�U�   �}�   um�E�Pj �M�����P�MQ�UR��,���P�MQ���������@�U�E�M�Q�UR�EP�MQ��D���R�EP�t�������P�M�U�E�    �5�E�Pj �M��D���P�MQ�UR��4���P�MQ�[�������@�U�E�M0+M�Q�U�R�M��
���P�EP�MQ��L���R�EP�!�������P�M�Uj j �M�e����E�P�MQ�UR�EP�MQ�UR��������E��M������E������M�������E�M�d�    Y[�M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �x���E�h  h���M�Qj��������E��E�    �}� t:j �M�_	��P�M�������E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]��������������������������������������������������������������������������U��j�h$�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �8���E�hD  h���M�Qj�������E��E�    �}� t:j �M���P�M������E��U��U��E��E����E��M�Q�M��?����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h�   h���M�Qj�_������E��E�    �}� t<jj �M����P�M��s����E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]������������������������������������������������������������������������U���`���3ŉE�VW�M̍E�P������   ���}��   �uЋ}�E_^�M�3��0�����]� ���������������������������������U��Q�M������]�����������������U��j�h��d�    P��   ���3ŉE�VP�E�d�    �M����% 0  = 0  u%�EP�MQ�UR�EP�MQ�UR��������  ��\���P�M�>�����l�����l�����d����E�    ��d���R�������E��E�������\���������E�P�M��0���E�   �M�M��E� ��`���R�M�������h�����h�����p����E���p���Q�I�������x����E���`��������U�R�   k���D�Q�   k� D�P��x��������MQ�UR�����������t�h�M�[����Ⱥ   k��T�;�u�E�� +�M����M��M�����3�M�&����и   k�
�D�;�u�M��-�U����U��M�~����E� �E�    �E�    j �M��G����E��E����t�U������   ��E��M�8����MQ�UR�)���������te�M������Q�U�R��������E��}�
sD�}�$|�E����E��.�}� u�}� u� �M��U���D���M����M��U����U��x����  �M��c�����u�E� ��M������E��E��E�j j�M�������E��E�    ��M�s����MQ�UR�d�����������   �M�������Q�U�R��������E��}�
s~�E��}�$|�E����E��.�}� u�}� u� �M��U���D���M����M��U����U��E�P�M��j������t%�U�R�M��V�����|�����|��������|����
�G�E�P�M��/������t�U���t�M�������M�;�t��j j�M��S����U����U�������}� u�"�E�P�M���������~�U����U���E��E���u�}� vy�M����u�l�e�E����E�t�M��1�U�R�M������ ;�u�}� u�M��1�U�R�M��l���� ;�}�E���   �� �U��
��~	�M����M��y����E��M������U���t�}� u�E�� 0�M����M��UR�EP�������ȅ�tB�M��������M��������;�u(�-����   k� � �M����E����E��M�:����}� uj��E��M�&����MQ�UR����������t'�M�����Ⱥ   k� �T�;�u�E����E�붃}� }�M��0�U����U��E����E���E��M�����MQ�UR����������tI�M������Q�U�R�K������E��}�
s(�}�$} �E��M���D���E����E��M����M���U�����  �EP�MQ�A������Ѕ���  �M�������   k��L�;�t �M�����и   k��D�;��i  �M��e�U����U��M������E� �E�    �EP�MQ�������Ѕ�t�h�M�3������   k��L�;�u�U��+�E����E��M�����3�M������Ⱥ   k�
�T�;�u�E�� -�M����M��M�V����UR�EP�G������ȅ�t*�M�����и   k� �D�;�u�E��M������M���t�U��0�E����E���E��M������MQ�UR�����������tI�M�N�����Q�U�R�������E��}�
s(�}�} �E��M���D���E����E��M����M���U���u�E���u�M�M��U�� �E���t����E������M��7�����t����M�d�    Y^�M�3��������]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hf�d�    P��   ���3ŉE�VP�E�d�    ��P���P�M�g�����`�����`�����X����E�    ��X���R�������t����E�������P��������E�P��t����S����E�   ��T���Q�M������\�����\�����d����E���d���P�v�������l����E���T��������M�Q�   k���P�   k� �¬�R��l��������E�E��E� �MQ�UR�����������t�h�M�~����Ⱥ   k��T�;�u�E�� +�M����M��M������3�M�I����и   k��D�;�u�M��-�U����U��M�����E�� 0�M����M��U��x�E����E��E� �E�    ǅ|���    �MQ�UR�:���������u�M������Ⱥ   k� �T�;�t�b�EP�M�-���P�%������ȅ�tB�M�����и   k��D�;�t�M�v����Ⱥ   k��T�;�u
�M�������E�j �M�������x�����x������t��x��������   ��E��M�����MQ�UR����������tk�M�������Q�U�R�)������E��}�sJ�}�$|��|�������|����.�}� u�}� u� �M��U�������M����M��U����U��r����.  �M�������u�E� ���t��������E��E��E�j j�M��N����E��E�    ��M������MQ�UR������������   �M�&�����Q�U�R�W������E��}���   �E��}�$|��|�������|����.�}� u�}� u� �M��U�������M����M��U����U��E�P�M��������t%�U�R�M�������p�����p��������p����
�G�E�P�M��~������t�U���t�M�b������M�;�t��j j�M������U����U�������}� u�"�E�P�M��*������~�U����U���E��E�����   �}� ��   ��x������u�{�t�E����E�t��x����1�U�R�M������� ;�u"�}� u"��x����1�U�R�M������ ;�}�E��%�   �� ��x����
��~��x�������x����_����E��M�������U���t�}� u�E�� 0�M����M��UR�EP�������ȅ�tE�M�&�������t���������;�u(�_����   k� � �M����E����E��M�l����}� uy��E��M�X����MQ�UR�I���������t-�M�����Ⱥ   k� �T�;�u��|�������|���밃�|��� }�M��0�U����U���|�������|�����E��M������MQ�UR�����������tI�M�=�����Q�U�R�n������E��}�s(�}�$} �E��M�������E����E��M����M���U�����  �EP�MQ�d������Ѕ���  �M��������   k��L�;�t �M�����и   k��D�;��i  �M��p�U����U��M�����E� �E�    �EP�MQ��������Ѕ�t�h�M�V������   k��L�;�u�U��+�E����E��M�����3�M�!����Ⱥ   k��T�;�u�E�� -�M����M��M�y����UR�EP�j������ȅ�t*�M������и   k� �D�;�u�E��M�:�����M���t�U��0�E����E���E��M�����MQ�UR����������tI�M�q�����Q�U�R�������E��}�s(�}�} �E��M�������E����E��M����M���U���u�E���u�M�M��U�� �E��|����ǅh���    �E������M��N�����h����M�d�    Y^�M�3��������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��   ���3ŉE�VP�E�d�    �EP�������x����M�Q��x����p����E�    �M��j�����u�E� ���x��������E��U��U��EP��������X����M�Q�   k�$�P�   k� ��$�R��X���������E�E��MQ�UR� ���������t�h�M�����Ⱥ   k��T�;�u�E�� +�M����M��M�����3�M�{����и   k��D�;�u�M��-�U����U��M�ӿ���E%   �E�}   u	�E�   �F�}   uǅd���   �(�} uǅl���    �
ǅl���
   ��l�����d�����d����U��E��E��E� �E� �MQ�UR�S�����������   �M�����Ⱥ   k� �T�;���   �E��M�����EP�MQ�������Ѕ�tY�M�y������   k��L�;�t�M�]����и   k��D�;�u!�}� t�}�u�E�   �E� �M譾����}� u�E�   �}� t0�}�
t*�}�uǅt���   �
ǅt���   ��t�����h����
ǅh���
   ��h�����`����E�Pj�M������E��E�    �   k�U��\�����M�����EP�MQ�������Ѕ���   �M�w�����P�M�Q��������p�����p���;�`���sz�E���p�����$���E���u�M����0t�E�;�\���s�M����M��E��E��U�R�M������ ��t$�M�Q�M��������|�����|������|�����G�U�R�M��ҽ��� ��t�M���t�M�������E�;�t��j j�M�������M����M�������}� u�"�U�R�M��~���� ��~�M����M���E� j �M�������E��U���t�}� vy�E����u�l�e�U����U�t�E��0�M�Q�M��!����;�u�}� u�E��0�M�Q�M������;�}�E� ��   �� �M����~	�E����E��y����M���t�U���u�E�� 0�M����M���U���u�E�E��M�� �U���T����E� �M�������E������M��������T����M�d�    Y^�M�3�������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M��F�����]�����������������U��Q�M��M���,�,�����]�����������U��Q�M�� ���]�����������������U����E�E��M��%�U����U��E�� t�M��+�U����U��E��t�M��#�U����U��   k� �U�
��Lt�   k� �E��M���E����E��-�M��I�U����U��E�� 6�M����M��U��4�E����E��M��   �M�}�   u�E�o�:�}�   t�   �� �E��M���U��t�E�X��E�x�E��E��M��M��U��E���M����M��U�� �E��]��������������������������������������������������������������������������������������U����M��E��8 t,�M��	�����E������E�U�R�E�P��������ȅ�t�U��    �E��@��M��A ��]�����������������������U��Q�M���]� ���U��Q�M���]� ���U��j�h �d�    PQ��   ���3ŉE�SVWP�E�d�    �e��M��M������E��E�P�M������M��A    �U��B    �E��@    �E�    �M��t	�E��Q�	�U��B�E��M�Q�M�}�����p�����p���Rj �E�P�1�������x����M���x����Q�M������E��E�Pj �M�Q��������|����U���|����B�M臶����t����M�Qj ��t���R�ͼ�����E��E��M��H��M�����j j �������u��E�������E������U��t.�E�Pj j.��������M��A�U�Rj j,�޶�����M��A���,�   �u����U�Rj �M��	����M�d�    Y_^[�M�3�������]� ��������������������������������������������������������������������������������������������������������������������U��j�h`�d�    P��   ���3ŉE�P�E�d�    h�  h���EP�������}$ v�M ���+t�E ���-u	�E�   ��E�    �U��U��M�R���%   =   u@�E���;E$w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M��U�R�M������|�����|�����t����E�    ��t���Q� ������E��E������M��E���j �U$R�M��D����E�   j �M��H���P�E E$P�   k� U R�M��<����E�P�M������x�����x����M��E��U�R�������E��E��M��Щ���E�P�M������E�j �M��;����E��M����ty�E����~o�M��L����E��U����tY�M����~O�E���U$+U�;�s?�E���U$+щU$�E�Pj�M$Q�M�������   �� �E����~	�U����U�뜍M��{����E$�M������E��U��}� |%�}� v�M�����;E$v�M�����+E$�E���E�    �E��E��M�Q���%�  �E��}�@ty�}�   tp�M�Q�UR�EP�MQ��T���R�EP�˲������P�M�U�E�    �E�Pj �M�蝳��P�MQ�UR��l���P�MQ贫������@�U�E�   �}�   um�M�Qj �M��Z���P�UR�EP��D���Q�UR�q�������P�M�U�E�P�MQ�UR�EP��\���Q�UR��������P�M�U�E�    �5�E�Pj �M�����P�MQ�UR��L���P�MQ��������@�U�E�M$+M�Q�U�R�M�賲��P�EP�MQ��d���R�EP�ʪ������P�M�Uj j �M�����E�P�MQ�UR�EP�MQ�UR�m������E��M�謸���E������M�蝸���E�M�d�    Y�M�3��Q�����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P�����3�P�E�d�    j �M�苵���E�    �E�(   �E�H;M��   �U���U��}�(s�E�(   h�   hȂj�E���P�M�QR�۽�����E�}� u�o����E�M�H��U�B���M�A�U�B;E�s�M�Q�E�H��    �ыU��M�P�ҋE�H�U�<� t(�E�H�U���M�Q�M� ���P��P�N������E�H�U�E���E������M�������M�d�    Y��]������������������������������������������������������������������������������������U��j�h��d�    P��D���3�P�E�d�    �E;��u<h8p�M������E�    j �MQj?�U�R�������E������M�������   j �M�贳���E�   �E�x v}jhhȂj�M�Q��R�`������E�E�M�H�}� u蹲���U�B�E��}� v<�M����M��U�B�M����U�E�H�U��E���}� t�M��M�B����E������M��j����M�d�    Y��]��������������������������������������������������������������������������������U����E�    �} u
hTQ������   k� �U�
��*u�   �� �U�
��u�|�} uj j �$������E��e�}?u�MQj �������E��L�E�    �	�U����U��}�#�   �M�����#Et�MQ�U�R��������΋EPj �������E��}� uh4p�M��,�����,h4p�M��,脷��P���������t�M�Q�M��,�����E��]��������������������������������������������������������������������U���j j �������E��}� u	�E��Q��E��E��M�Q�M��$�^����UR�EP�MQ��������]��������������������������������U��j�h��d�    P��P���3�P�E�d�    j j ��������   ������#Uu�   �} um�����E�jJhȂ�E�Pj�������E��E�    �}� tj �MQ�M�蠺���E���E�    �U�U��E��������膬��P�E�P�M�~���� ����m���P�MQ������P�M�\���j j �������   ������#Uu�   �} um������E�jKhȂ�E�Pj�d������E��E�   �}� tj �MQ�M������E���E�    �U�U��E������\��ҫ��P�E�P�M�ʺ��� �\�蹫��P�MQ������P�M診��j j �5������   ������#Uu�   �} um�F����E�jLhȂ�E�Pj谲�����E��E�   �}� tj �MQ�M��w����E���E�    �U܉U��E������`�����P�E�P�M����� �`�����P�MQ�%�����P�M�����j j �N������   ������#Uu�   �} uo�����E�jMhȂ�E�Pj��������E��E�   �}� tj j �MQ�M������E���E�    �UԉU��E���������h���P�E�P�M�`���� ����O���P�MQ������P�M�>���j j �������   ������#Uu�   �} um������E�jOhȂ�E�Pj�F������E��E�   �}� tj �MQ�M�������E���E�    �ỦU��E��������贩��P�E�P�M謸��� ���蛩��P�MQ蕾����P�M芸���UR�EP�MQ�UR�������EP�MQ�UR�EP�[������MQ�UR�EP�MQ��������U�BE�M�A�M����P�M�������E�M�d�    Y��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��E��8 t,�M��	�����E������E�U�R�E�P��������ȅ�t�U��    ��E�P��������M��A�U��B�E��@��]��������������������������������������U����E���E�M�����M���M�} v�U�P�M�����������ȋM�U��E�A�E]���������������������������������U����E���E�M蠚���} v�MQ�M�������3����ӋU�E��M�J�E]����������������������������U��Q�M��E��8 tj�M��R葬�����E��     ��]���������������������U��Q�M��E��HQ�W������U��BP�H������M��QR�9�������]�������������������������U����M��E�;Eu�a�M�Q�M����P�U�R�M�����P蚻��������t�M�yr�UR�M�������!j j�M��]����EP�������P�M������E���]� �����������������������������������U��Q�M��@QPj �MQ�M�������]� ���������������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E��@��]����������������U����M��E�    �E��HQ�M�~����U����U��E��]� ���������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP�4������E�    �M�Q�M�b����E��U��U��E�    �E�P�M����P�MQ�UR�E�P�M�Q�0������E��E������M������   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R�������E̍EP�MQ�6������Ѕ�t�E ����U �
�E�;E�t�}� u	�}���  v�M ����E ��,�   k� �DЃ�-u
3�+M̉M���ỦUċE$f�M�f��U�E��M�J�E�M�d�    Y�M�3��u�����]�  ������������������������������������������������������������������������������������������������������U��j�h�d�    P��P���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP�D������E�    �M�Q�M�r����E��U��U��E�    �E�P�M�����P�MQ�UR�E�P�M�Q�@������E��E������M������   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R�������E̍EP�MQ�F������Ѕ�t�E ����U �
�E�;E�t�}� u�}��v�M ����E ��*�   k� �DЃ�-u
3�+M̉M���ỦUċE$�Mĉ�U�E��M�J�E�M�d�    Y�M�3�芷����]�  �����������������������������������������������������������������������������������������������������������U��j�hX�d�    P��@���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP�T������E�    �M�Q�U�R�M�~����E��E��E��E�    �M�Q�M�����P�UR�EP�M�Q�U�R�L�����P�E�P�M�Q�������E��E������M������UR�EP肻�����ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3�������]�  �������������������������������������������������������������������������������U��j�h��d�    P��@���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP��������E�    �M�Q�U�R�M������E��E��E��E�    �M�Q�M�M���P�UR�EP�M�Q�U�R�̛����P�E�P�M�Q�\������E��E������M�薒���UR�EP�������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3��n�����]�  �������������������������������������������������������������������������������U���T���3ŉE��M�h)  h���EP�MQ�UR�EP�l������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q�&�����P�U�R�E�P赶�����]��}� t�M���QQ�E��$謹�����]��UR�EP褸�����ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3�������]�  ����������������������������������������������������������������������������U���X���3ŉE��M�hA  h���EP�MQ�UR�EP�������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q�֪����P�U�R�E�P�L������]��}� t�M���Q���E��$趎�����]��UR�EP�R������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��ɱ����]�  ��������������������������������������������������������������������������U���X���3ŉE��M�hY  h���EP�MQ�UR�EP��������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q膩����P�U�R�E�P�Q������]��}� t�M���Q���E��$�F������]��UR�EP�������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��y�����]�  ��������������������������������������������������������������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�hq  h���EP�MQ�UR�EP�d������E�    �M�Q�M蒴���E��U��U��E�    �E�Ph   �MQ�UR�E�P�M�Q�d������E��E������M��?����   ��t"�E�P�M�Q�U�R�E�P�ҽ����3ɉE��M���U�R�E�P�M�Q�U�R�p������E��U��E��E��M��M��UR�EP�V������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E��M$��U�E��M�J�E�M�d�    Y�M�3��®����]�  ���������������������������������������������������������������������������������������������������U��j�h�d�    P��D���3ŉE�P�E�d�    �M�h   h���EP�MQ�UR�EP�������E�    �M�Q�U�R�M農���E��E��E��E�    �M�Q�M����P�UR�EP�M�Q�U�R茔����P�E�P�M�Q�&������E��U��E������M��S����UR�EP迲�����ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3��%�����]�  ��������������������������������������������������������������������������������������U��j�hX�d�    P��D���3ŉE�P�E�d�    �M�h  h���EP�MQ�UR�EP�������E�    �M�Q�U�R�M�.����E��E��E��E�    �M�Q�M�}���P�UR�EP�M�Q�U�R�������P�E�P�M�Q�L������E��U��E������M��É���UR�EP�/������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3�蕫����]�  ��������������������������������������������������������������������������������������U��j�h��d�    P��   ���3ŉE�P�E�d�    ��L���h�  h���EP�MQ�UR�EP�n�����ǅx��������M����% @  �'  ��H���Q�M胯����\�����\�����P����E�    ��P���P�#�������p����E�������H����3���j j�M��4����E�   ��|���Q��p����������@�����@�����8����E���8���P�M��E����E���|����U���j �M��t����M�Q��p���������d�����d�����<����E���<���P�M�������E��M������M�����Pj�MQ�UR�Z�������x����E������M��ۘ���   ǅh���    ��h���P��`���Q�M�K�����T�����T�����D����E�   ��D���P�M����P�MQ�UR�E�P��L���Q�
�����P��X���R�E�P藷������l����E�������`����ˆ���M�9�X���t��h��� u��l���w��l�����x����EP�MQ�������Ѕ�t�E ����U �
��x��� }�E ����U �
�*��x��� tǅt���   �
ǅt���    �E$��t�����U�E��M�J�E�M�d�    Y�M�3��]�����]�  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��E�    �E��HQ�M������U����U��E��]� ���������������U���P���3ŉE��M��EP�M�n���Ph��M�Q�U�R�φ����Pj@�E�P������P�M�Q�UR�EP�MQ�UR�EP�M�Q触���� �E�M�3�������]� �����������������������������������U���P���3ŉE��M��EP�M�����Ph��M�Q�U�R�/�����Pj@�E�P�������P�M�Q�UR�EP�MQ�UR�EP�M�Q������ �E�M�3��B�����]� �����������������������������������U���   ���3ŉE���`����M������T�����X�����X��� 0|	��T��� w%�M����%    uǅh���   ǅl���    ��M�������h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M�P���% 0  =    �  �E��^�E������D��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E�(�����u��x����  s�E�5��]���E�x^����Aud���t�����
��t����}� |M	��|���
rB���]����u2��t����  s&�E���]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M����Pj �E�P��`���Q讂����Pjl�U�R�&�����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P�������,�E�M�3��q�����]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE���`����M������T�����X�����X��� 0|	��T��� w%�M����%    uǅh���   ǅl���    ��M�o�����h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M�����% 0  =    ��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E�(�����u��x����  s�E�5��]���E�x^����Aud���t�����
��t����}� |M	��|���
rB���]����u2��t����  s&�E���]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M�����PjL�E�P��`���Q�g����Pjl�U�R�߻����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P趍����,�E�M�3��*�����]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���H���3ŉE��M��EPh �j@�M�Q蹺����P�U�R�EP�MQ�UR�EP�MQ�U�R������ �E�M�3�������]� �����������������������������U���P���3ŉE��M��E P�MQ�M�
���Ph��U�R�E�P�k~����Pj@�M�Q������P�U�R�EP�MQ�UR�EP�MQ�U�R�C����� �E�M�3��~�����]� �����������������������������������������������U���P���3ŉE��M��E P�MQ�M�Z���Ph��U�R�E�P�}����Pj@�M�Q�k�����P�U�R�EP�MQ�UR�EP�MQ�U�R蓝���� �E�M�3��Ν����]� �����������������������������������������������U��j�h�d�    P��   ���3ŉE�VP�E�d�    �M�h�  h���EP�������M����% @  u4�MQ�UR�EP�MQ�UR�EP�M���M��B$�ЋE��  ��  ��p���Q�M�ˡ���E��U���|����E�    ��|���P�q������E��E�������p����z���M�������E�   �M��t%�U�R�M��.����E��E�P�M��Ӏ���M��ŋ���#�M�Q�M��#����E��U�R�M�讀���M�蠋���M�������t�����x�����x��� |:	��t��� v/�M�̧�����M��?���;�v�M趧�����M��)���+��u���E�    �E��E��M�4���%�  ��@t6�M�Q�UR�EP�MQ��`���R�E�P軃������P�M�U�E�    �M��Ŏ��P�M��Є��P�EP�MQ��h���R�E�P�|������P�M�Uj j �M�����E�P�MQ�UR�EP�MQ�U�R�D������E������M�耊���E�M�d�    Y^�M�3��3�����]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M��E��@��]����������������U����M��E�    �E��HQ�M讽���U����U��E��]� ���������������U����M��E��H��u�M��<����U�B��u�M�)����M��9 u�U�: t�E��8 t�M�9 u	�E�    ��E�   �E���]� ����������������������������������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�P�M��t���P�M�-����E��]� ���������U��j�h`�d�    P�����3�P�E�d�    �E�    �M��F����E�    j �M��e����E������E��E�M�;��   �U���M��P��P�ي�����E��M��U�R�Ǘ�����E���M��B�ЋM��Q��?�U�}�?u�M���請��Pj 讲�����C�E�    �	�E���E�}�+�   �M�����#U�t�M����j���P�E�P�k������ƍM�Q�M�5����U����U��E� �M��ذ���E������M��u���E��E������M��u���M�d�    Y��]�������������������������������������������������������������������������������������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E��H;Ms�M������U��@Q+B;Ew�M��&����} vo�M��QU�U�j �E�P�M��W���ȅ�tN�U��B+EP�M��K���EP�M��?���EEP�7������MQ�UR�EP�M��r���M�Q�M�����E���]� ����������������������������������������������U��Q�M��M��A�Q��]�������������U����M��M��y����E�U��}� |,�}� v$�M������E��E��M��U�R臶�����E���EP�v�����P�M���M��B�ЉE�E��]� ���������������������������������U��Q�M��E���M��B�Ћ�]���������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��EP�MQ�UR�E���M��B�Ћ�]� ����������U����M��E��H �M�P$�U��E��M�H �U�P$�E�U���]� �������������U��Q�M��M��A �Q$��]�������������U��Q�EP�E���$�&q�����]��E���]��������������U��EP���E�$��p����]�������U���8���3ŉE�VW�E�    3��EԉE؉E܉E��E�E�E�E��E�E������E��m����E���u���   ��< u	�E�   ��E�    �UȉU؃}� uQ�E�    �	�Ẽ��É}�   }6�M�Q�ڂ������t$�U����M̃��   ���L�ȋU����L�븹   �uЋ}�E_^�M�3�腓����]�������������������������������������������������������������������������U���d���3ŉE�VW�E�x t0�M���   ~蕺��� *   ����   �U�E��   �t�r�E�    �} u�M�Q�������   ���}��UЉU�E�Pj �M�QR�EPj�MQj �U�P� �Ẽ}� t�}� t����� *   �����E�_^�M�3��p�����]����������������������������������������������������U��EP�MQ�UR�EP�d�����]�������������������U��]����������U��EP�M�N���]����������������U��Q�EP�M��T���P�MQ�M��G���P��������]�����������������������U��Q�EP�M�����P�MQ�M�����P�O�������]�����������������������U��EP�M�K���]����������������U��]����������U��Q�EP�MQ�g������Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ�K������Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ��}�����Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ赍�����Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ�x�����Ѕ�u	�E�   ��E�    �E���]���������������U��Q�EP�MQ豎�����Ѕ�u	�E�   ��E�    �E���]���������������U��Q�E�    �} u�%�}���w�E��P�Å�����E��}� u�9|���E���]������������������U��Q�E�    �} u�%�}���w�E��P�s������E��}� u��{���E���]������������������U��Q�EP�MQ�v�����E��U�R�EP�MQ�UR�EP�MQ�������E��]������������������U��Q�EP�M�Q��w�����UR�E�P�-m�����M�Q�U�R�EP�MQ�UR�EP�MQ�׺�����E��]��������������������������������U����M臶���E���E�M;Mt�U�P�M�������茞���ϋM�U��E�A�E]������������������������U��EP�MQ�UR�EP�MQ�M������E]�������������U��Q�EP�MQ��k�����E��U�R�EP�MQ�UR�EP�MQ�������E��]������������������U��Q�EP�M�Q�pp�����UR�E�P��k�����M�Q�U�R�EP�MQ�UR�EP�MQ�������E��]��������������������������������U����M�ex���E���E�M;Mt�U�P�M�������Ø���ϋM�U��E�A�E]������������������������U��EP�MQ�UR�EP�MQ�L������E]�������������U��} u�EP�MQhH]�V����]�����������������U��} u�EP�MQhH]�&����]�����������������U��} u�EP�MQhH]��~����]�����������������U��} u�EP�MQhH]��~����]�����������������U��} u�EP�MQhH]�~����]�����������������U��]������������U��]������������U��} u�EP�MQhH]�F~����]�����������������U��} u�EP�MQhH]�~����]�����������������U��E;EtE�MQ�UR�EP�������MQ�UR�EP�٧�����M;Ms�UR�EPh�]�}����]�������������������������������U��E;EtE�MQ�UR�EP�������MQ�UR�EP�������M;Ms�UR�EPh�]�D}����]�������������������������������U��E;EtE�MQ�UR�EP赐�����MQ�UR�EP衐�����M;Ms�UR�EPh�]��|����]�������������������������������U��E;EtE�MQ�UR�EP蔑�����MQ�UR�EP耑�����M;Ms�UR�EPh�]�d|����]�������������������������������U��E;EtE�MQ�UR�EP聎�����MQ�UR�EP�m������M;Ms�UR�EPh�]��{����]�������������������������������U��Q�EP�MQ�+������E��U��U���]����������������U��Q�EP�MQ�q�����E��U��U���]����������������U��Q�EP�M�Q膑�������P�MQ�UR�EP�MQ�ev������]���������������������������U��Q�EP�M�Q����������P�MQ�UR�EP�MQ�A�������]���������������������������U��Q�EP�M�Q�Mf�������P�MQ�UR�EP�MQ��������]���������������������������U��Q�EP�M�Q�p�������P�MQ�UR�EP�MQ��������]���������������������������U��Q�EP�M�Q�t�������P�MQ�UR�EP�MQ��y������]���������������������������U��Q�EP�k�����E��M�Q�UR�EP�MQ�UR�EP�MQ蘵������]���������������������U��Q�EP��m�����E��M�Q�UR�EP�MQ�UR�EP�MQ�z������]���������������������U��Q�E�E��	�M����M��U����t�M���E;�t�݋E�+E����]����������������������U��Q�E�E��	�M����M��U����t�M���E;�t�݋E�+E����]����������������������U��j�h��d�    P��D���3ŉE�VP�E�d�    �E�    �	�E����E��MM����t'�EE���   k� �U�;�u	�M���M��j �UR�M���x���E�    �E������E�   ��Eă��EċM衑���E������E� �E�    �E�    �	�Mȃ��MȋU�;U�#  �	�EЃ��EЋMM����t�EE���   k� �U�;�t�̋M�Q�M��]m�����t�E�P�M��Jm���MЉM��   �U�UĉUЋEE���   k� �U�;�t�MM����u.�}�s�EĉE���E�   �M�Q�M���l���U���EȉE��[�MQ�UR�g���������u�MM��1�M��}����;�t(�}�s�EĉE���E�   �M�Q�M��l���U����E�������Eυ�t�MQ�UR�����������t��v����M��M��E������M��r���E��M�d�    Y^�M�3��M�����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��D���3ŉE�VP�E�d�    �E�    �	�E����E��MM����t'�EE���   k� �U�;�u	�M���M��j �UR�M���u���E�    �E������E�   ��Eă��EċM�����E������E� �E�    �E�    �	�Mȃ��MȋU�;U�#  �	�EЃ��EЋMM����t�EE���   k� �U�;�t�̋M�Q�M��mj�����t�E�P�M��Zj���MЉM��   �U�UĉUЋEE���   k� �U�;�t�MM����u.�}�s�EĉE���E�   �M�Q�M���i���U���EȉE��[�MQ�UR�i��������u�MM��1�M������;�t(�}�s�EĉE���E�   �M�Q�M��i���U����E�������Eυ�t�MQ�UR�i��������t��v����M��M��E������M��o���E��M�d�    Y^�M�3��]�����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��D���3ŉE�VP�E�d�    �E�    �	�E����E��M��U�J��t(�M��U�J�   k� �M�;�u	�E���E��j �MQ�M�� s���E�    �E������E�   ��Uă��UċM迋���E������E� �E�    �E�    �	�Eȃ��EȋM�;M�(  �	�UЃ��UЋEЋM�A��t�EЋM�A�   k� �E�;�t�ʋU�R�M��yg��� ��t�M�Q�M��fg���UЉU��   �E�EĉEЋMЋU�J�   k� �M�;�t�EЋM�A��u.�}�s�EĉE���E�   �M�Q�M��g���U���EȉE��\�MQ�UR聃��������u�MЋU�4J�M�x����;�t(�}�s�MĉM���E�   �U�R�M��f���M����E�������Uυ�t�EP�MQ�������Ѕ�t��q����E��E��E������M��l���E��M�d�    Y^�M�3��f}����]����������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hX�d�    P��D���3ŉE�VP�E�d�    �E�    �	�E����E��M��U�J��t(�M��U�J�   k� �M�;�u	�E���E��j �MQ�M��p���E�    �E������E�   ��Uă��UċM�����E������E� �E�    �E�    �	�Eȃ��EȋM�;M�(  �	�UЃ��UЋEЋM�A��t�EЋM�A�   k� �E�;�t�ʋU�R�M��d��� ��t�M�Q�M��vd���UЉU��   �E�EĉEЋMЋU�J�   k� �M�;�t�EЋM�A��u.�}�s�EĉE���E�   �M�Q�M��d���U���EȉE��\�MQ�UR�c��������u�MЋU�4J�M�&�����;�t(�}�s�MĉM���E�   �U�R�M��c���M����E�������Uυ�t�EP�MQ�1c�����Ѕ�t��q����E��E��E������M���i���E��M�d�    Y^�M�3��vz����]����������������������������������������������������������������������������������������������������������������������������������������������������������U����M��E��H(��t�U�B�E��	�M�Q�U��E���,Pj �M�Q�Y�����U��B�E�H.��v	�E��Q�	�U�B �E�M���,Qj �U�R�cY�����M��A�U�B/��v	�E��	�M�Q$�U��E���,Pj �M�Q�*Y�����U��B�E���,Pj �   k� �E�H�R�Hu�����M�f�A�U���,Rj �   k� �U�B�Q�u�����U�f�B��]� �������������������������������������������������������������������������������U��Q�M��EPj �   k� �E��R�t�����M�f�A�URj �   k� �U�B�Q�rt�����U�f�B��]�4 ������������������������������������U���4���3ŉE�VW�M̍E�P�M�#����}̃��   ���M̃�Qj �M�Y��P�W�����ỦB�Ẽ�Pj �M�V��P�W�����M̉A�Ũ�Rj h���sW�����M̉A_^�M�3��aw����]� ��������������������������������������������������U����M��E��H(��t�U�B8�E��	�M�Q<�U��E�P�5S�����M��A�U�B.��v	�E����	�M�QH�U�E�P�S�����M��A�U�B/��v	�E��	�M�QL�U��E�P��R�����M��A�   k� �M�Q@�M�f�f�Q�   k� �U�BD�U�f�f�B��]� ��������������������������������������������������������������U��Q�M��   k� �U�B0�U�f�f�B�   k� �E�H4�E�f�
f�H��]�4 �����������������U���4���3ŉE�VW�M̍E�P�M�����}̃��   ���M�W���P��Q�����M̉A�M�b��P�Q�����ỦBh��Q�����M̉A_^�M�3��Lu����]� ���������������������������������������������U��Q3��E��E���]�����������������U��Q3��E��E���]�����������������U��Q�E�M���E��]��������������U��Q�E�M���E��]��������������U��Q�E�M���E��]��������������U��Q�E�M���E��]��������������U��Q�E�M���E��]��������������U��Q�E���]������U��Q�E���]������U��E]���������U��E]���������U�����E���E�M���M�U;Ut8�E;Et0�M��E�;�}����M��U��M�;�}�   �4뮋E;Et	�E�������M;Mt	�E�   ��E�    �U��U��E���]�������������������������������������������������U��EP�MQ�UR�EP�MQ�X�����]����������������U��Q�E+E���E��M+M��9M�w!�U���R�EP�M+M����Q�UR� `�����E���]�����������������������������U��EP�MQ�UR�EP�MQ蕜����]����������������U���3�f�E��E�    �MQ�U�Rj�EP�M�Q�k�����f�E���]����������������������������U���3�f�E��E�    �MQ�U�Rj�EP�M�Q������f�E���]����������������������������U���,�E�    �EP�&}�������E�M�M��E�    �U�U���E�+E�E��M�M�M�U����U��}� v)�EP�M�Q�U�R�E�P�M�Q臠�����E�}� �붋U����U�h  h��Ɇ��P3ɋE��   �������Q�wP�����E؋E؉E��M��M��E�    �$�U�+U�U��EE�E�M����M��U���U�}� v)�EP�M�Q�U�R�EP�M�Q�������E�}� ��3ҋE�f��E���]������������������������������������������������������������������������������������U���,�E�    �EP�{�������E�M�M��E�    �U�U���E�+E�E��M�M�M�U����U��}� v)�EP�M�Q�U�R�E�P�M�Q�������E�}� �붋U����U�h�  h��I���P3ɋE��   �������Q��N�����E؋E؉E��M��M��E�    �$�U�+U�U��EE�E�M����M��U���U�}� v)�EP�M�Q�U�R�EP�M�Q�g������E�}� ��3ҋE�f��E���]������������������������������������������������������������������������������������U��Q�E���]������U��Q�E���]������U��E]���������U��E]���������U��E]���������U��j�h��d�    P��`���3�P�E�d�    �M��E�   ���̉eȍEP�`���E�M�M��E����̉e��UR�p`���E�E�E��E��M�Q�M��zQ���E�U�U��E����̉e��E�P�����E܋M܉M��E��U�R�M���_���E؋E؉E��E����̉e��U�R跛���E��E��M�迉���EЋEЉE��E��M��S���E��M��S���E� �M�S���E������M�xS���E̋M�d�    Y��]� �������������������������������������������������������������������������������������U��j�h8�d�    P��`���3�P�E�d�    �M��E�   ���̉eȍEP�d����E�M�M��E����̉e��UR�F����E�E�E��E��M�Q�M��hZ���E�U�U��E����̉e��E�P�S���E܋M܉M��E��U�R�M��ߍ���E؋E؉E��E����̉e��U�R�QS���E��E��M���f���EЋEЉE��E��M��Z���E��M��tZ���E� �M�hZ���E������M�YZ���E̋M�d�    Y��]� �������������������������������������������������������������������������������������U��Q�M��EP�ވ����P�MQ�U�R�Ό������]� ����������������������U��j�h��d�    P�����3�P�E�d�    �M�EPj�/k�����E��E�    �}� t�MQ�_������U�� ��M��M���E�    �U�U��E������M�d�    Y��]� ������������������������������������������U��EP������P�MQ�M����]�������������������U��Q�M��EP������P�MQ�U�R��X������]� ����������������������U��j�h��d�    P�����3�P�E�d�    �M�EPj�j�����E��E�    �}� t�MQ薏�����U�� ��M��M���E�    �U�U��E������M�d�    Y��]� ������������������������������������������U��EP�)�����P�MQ�M�_��]�������������������U��Q�E;Eu�M�U��E�A�E�{�yhQ  h8��MQ�UR�)e����hR  h8��EP�'V�����MQ�UR� E�����E��E�P�MQ�UR�EP�r����P�MQ�	r����P�UR�l�����E��]���������������������������������������������������U��Q�E;Eu�M�U��E�A�E�{�yhQ  h8��MQ�UR�Yd����hR  h8��EP�ő�����MQ�UR�g�����E��E�P�MQ�UR�EP�Fq����P�MQ�9q����P�UR�f�����E��]���������������������������������������������������U��Q�M��EP�M�Q�G������]� �������������������U��Q�M���]� ���U��EP�M�IZ��]����������������U��Q�M��EP�M�Q�������]� �������������������U��Q�M���]� ���U��EP�M�O��]����������������U��E]���������U��E]���������U��E]���������U��E]���������U��j�h��d�    P��$���3�P�E�d�    j �M���S���E�    �(��E���P���E�M�Q�M�iw���E�}� t�n�}� t�U��U��`�EP�M�Q�Of�������uh|]�M��Y��hH=�U�R�Oz���.�E��E�M��(��U��U�E��M�B�ЋM�Q�ۄ�����U�U��E������M��~���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h(�d�    P��$���3�P�E�d�    j �M��R���E�    ����E����N���E�M�Q�M�)v���E�}� t�n�}� t�U��U��`�EP�M�Q�h�������uh|]�M���W��hH=�U�R�y���.�E��E�M�����U��U�E��M�B�ЋM�Q蛃�����U�U��E������M��W}���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hX�d�    P��$���3�P�E�d�    j �M��{Q���E�    ���E���M���E�M�Q�M��t���E�}� t�n�}� t�U��U��`�EP�M�Q��f�������uh|]�M��V��hH=�U�R��w���.�E��E�M����U��U�E��M�B�ЋM�Q�[������U�U��E������M��|���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��;P���E�    ����E���XL���E�M�Q�M�s���E�}� t�n�}� t�U��U��`�EP�M�Q��]�������uh|]�M��KU��hH=�U�R�v���.�E��E�M�����U��U�E��M�B�ЋM�Q�������U�U��E������M���z���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M���N���E�    ����E���K���E�M�Q�M�ir���E�}� t�n�}� t�U��U��`�EP�M�Q�:S�������uh|]�M��T��hH=�U�R�Ou���.�E��E�M�����U��U�E��M�B�ЋM�Q�������U�U��E������M��y���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��M���E�    ����E����I���E�M�Q�M�)q���E�}� t�n�}� t�U��U��`�EP�M�Q�]�������uh|]�M���R��hH=�U�R�t���.�E��E�M�����U��U�E��M�B�ЋM�Q�~�����U�U��E������M��Wx���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M��{L���E�    ���E���H���E�M�Q�M��o���E�}� t�n�}� t�U��U��`�EP�M�Q��}�������uh|]�M��Q��hH=�U�R��r���.�E��E�M����U��U�E��M�B�ЋM�Q�[}�����U�U��E������M��w���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hH�d�    P��$���3�P�E�d�    j �M��;K���E�    ����E���XG���E�M�Q�M�n���E�}� t�n�}� t�U��U��`�EP�M�Q�_�������uh|]�M��KP��hH=�U�R�q���.�E��E�M�����U��U�E��M�B�ЋM�Q�|�����U�U��E������M���u���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hx�d�    P��$���3�P�E�d�    j �M���I���E�    ���E���F���E�M�Q�M�im���E�}� t�n�}� t�U��U��`�EP�M�Q�?l�������uh|]�M��O��hH=�U�R�Op���.�E��E�M����U��U�E��M�B�ЋM�Q��z�����U�U��E������M��t���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��H���E�    ����E����D���E�M�Q�M�)l���E�}� t�n�}� t�U��U��`�EP�M�Q��6�������uh|]�M���M��hH=�U�R�o���.�E��E�M�����U��U�E��M�B�ЋM�Q�y�����U�U��E������M��Ws���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��{G���E�    ���E���C���E�M�Q�M��j���E�}� t�n�}� t�U��U��`�EP�M�Q�a�������uh|]�M��L��hH=�U�R��m���.�E��E�M����U��U�E��M�B�ЋM�Q�[x�����U�U��E������M��r���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M��;F���E�    ����E���XB���E�M�Q�M�i���E�}� t�n�}� t�U��U��`�EP�M�Q�96�������uh|]�M��KK��hH=�U�R�l���.�E��E�M�����U��U�E��M�B�ЋM�Q�w�����U�U��E������M���p���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h8�d�    P��$���3�P�E�d�    j �M���D���E�    ���E���A���E�M�Q�M�ih���E�}� t�n�}� t�U��U��`�EP�M�Q���������uh|]�M��J��hH=�U�R�Ok���.�E��E�M����U��U�E��M�B�ЋM�Q��u�����U�U��E������M��o���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hh�d�    P��$���3�P�E�d�    j �M��C���E�    ���E����?���E�M�Q�M�)g���E�}� t�n�}� t�U��U��`�EP�M�Q�Yp�������uh|]�M���H��hH=�U�R�j���.�E��E�M����U��U�E��M�B�ЋM�Q�t�����U�U��E������M��Wn���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��{B���E�    ����E���>���E�M�Q�M��e���E�}� t�n�}� t�U��U��`�EP�M�Q�S�������uh|]�M��G��hH=�U�R��h���.�E��E�M�����U��U�E��M�B�ЋM�Q�[s�����U�U��E������M��m���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��;A���E�    ����E���X=���E�M�Q�M�d���E�}� t�n�}� t�U��U��`�EP�M�Q�WJ�������uh|]�M��KF��hH=�U�R�g���.�E��E�M�����U��U�E��M�B�ЋM�Q�r�����U�U��E������M���k���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M���?���E�    ����E���<���E�M�Q�M�ic���E�}� t�n�}� t�U��U��`�EP�M�Q�a�������uh|]�M��E��hH=�U�R�Of���.�E��E�M�����U��U�E��M�B�ЋM�Q��p�����U�U��E������M��j���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h(�d�    P��$���3�P�E�d�    j �M��>���E�    ����E�x���:���E�M�Q�M�)b���E�}� t�n�}� t�U��U��`�EP�M�Q��o�������uh|]�M���C��hH=�U�R�e���.�E��E�M�����U��U�E��M�B�ЋM�Q�o�����U�U��E������M��Wi���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hX�d�    P��$���3�P�E�d�    j �M��{=���E�    � ��E���9���E�M�Q�M��`���E�}� t�n�}� t�U��U��`�EP�M�Q�#8�������uh|]�M��B��hH=�U�R��c���.�E��E�M�� ��U��U�E��M�B�ЋM�Q�[n�����U�U��E������M��h���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��;<���E�    ����E�|��X8���E�M�Q�M�_���E�}� t�n�}� t�U��U��`�EP�M�Q�/�������uh|]�M��KA��hH=�U�R�b���.�E��E�M�����U��U�E��M�B�ЋM�Q�m�����U�U��E������M���f���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M���:���E�    ���E����7���E�M�Q�M�i^���E�}� t�n�}� t�U��U��`�EP�M�Q�E�������uh|]�M��@��hH=�U�R�Oa���.�E��E�M����U��U�E��M�B�ЋM�Q��k�����U�U��E������M��e���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��9���E�    ����E�t���5���E�M�Q�M�)]���E�}� t�n�}� t�U��U��`�EP�M�Q�L�������uh|]�M���>��hH=�U�R�`���.�E��E�M�����U��U�E��M�B�ЋM�Q�j�����U�U��E������M��Wd���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M��{8���E�    � ��E���4���E�M�Q�M��[���E�}� t�n�}� t�U��U��`�EP�M�Q�+�������uh|]�M��=��hH=�U�R��^���.�E��E�M�� ��U��U�E��M�B�ЋM�Q�[i�����U�U��E������M��c���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hH�d�    P��$���3�P�E�d�    j �M��;7���E�    ����E���X3���E�M�Q�M�Z���E�}� t�n�}� t�U��U��`�EP�M�Q�NN�������uh|]�M��K<��hH=�U�R�]���.�E��E�M�����U��U�E��M�B�ЋM�Q�h�����U�U��E������M���a���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hx�d�    P��$���3�P�E�d�    j �M���5���E�    �$��E����2���E�M�Q�M�iY���E�}� t�n�}� t�U��U��`�EP�M�Q�+0�������uh|]�M��;��hH=�U�R�O\���.�E��E�M��$��U��U�E��M�B�ЋM�Q��f�����U�U��E������M��`���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��$���3�P�E�d�    j �M��4���E�    ����E�t���0���E�M�Q�M�)X���E�}� t�n�}� t�U��U��`�EP�M�Q��a�������uh|]�M���9��hH=�U�R�[���.�E��E�M�����U��U�E��M�B�ЋM�Q�e�����U�U��E������M��W_���E܋M�d�    Y��]��������������������������������������������������������������������������U��Q�M��EP�M��uP���E���]� ��������������������U��Q�M��M��e���E���]�����������U��Q�M��EP�M��%P���E���]� ��������������������U��Q�M��M��d���E���]�����������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��I���E�    �M�����U��E�B(�MQ�UR�M���:���E������E��M�d�    Y��]� �����������������������������������������U��j�h�d�    PQ���3�P�E�d�    �M��EP�M���H���E�    �M�����U��E�B(�MQ�UR�M��.���E������E��M�d�    Y��]� �����������������������������������������U��j�h8�d�    PQ���3�P�E�d�    �M��M��I���E�    �M��)h���E������E��M�d�    Y��]� ������������������������U��j�hh�d�    PQ���3�P�E�d�    �M��M��k���E�    �M��Ni���E������E��M�d�    Y��]� ������������������������U��Q�M��EP�M��IK���M��U�B�A�E���]� ������������������������U��j�h��d�    PQ���3�P�E�d�    �M��M��q���E�    �EP�M��_]���M��U�Q�E������E��M�d�    Y��]� ���������������������������U��Q�M��M��Rq���E��@    �E���]�����������������U��Q�M��EP�M���.���M��U�B�A�E���]� ������������������������U��j�h��d�    PQ���3�P�E�d�    �M��M���_���E�    �EP�M��o\���M��U�Q�E������E��M�d�    Y��]� ���������������������������U��Q�M��M��_���E��@    �E���]�����������������U��Q�M��EP�M��po���E���]� ��������������������U��Q�M��EP�MQ�M��[-���E���]� ����������������U��Q�M��EP�M��*(���E���]� ��������������������U��Q�M��EP�MQ�M���m���E���]� ����������������U��Q�M��M��V���E��@    �M��A    �E���]�����������������������U��Q�M��M��PV���E��@    �M��A    �E���]�����������������������U��Q�M��EP�M���n���E���]� ��������������������U��Q�M��M���L���E���]�����������U��Q�M��EP�M��OY���E���]� ��������������������U��Q�M��M���R���E���]�����������U��Q�M��E���]� ����������������U��Q�M��E���]�������������������U��Q�M��E���]� ����������������U��Q�M��E���]�������������������U����M��E�P�M���P�M��q��j j �M��hb���MQ�oa����P�M��;W���E���]� ������������������������U��j�h��d�    P�����3�P�E�d�    �M�E�P�M�Q�M�#�����b��P�M������E�    j j �M���a�����Rj �EP�M��_���E������E�M�d�    Y��]� �������������������������������������U��j�h(�d�    P�����3�P�E�d�    �M�M���J��P�M��F���E�    j j �M��6a���EP�MQ�M��&���E������E�M�d�    Y��]� ����������������������������������������U��j�hX�d�    P�����3�P�E�d�    �M�M��2J��P�M�����E�    j j �M��`���EP�M��j���E������E�M�d�    Y��]� �����������������������������U��j�h��d�    P�����3�P�E�d�    �M�M��I��P�M�����E�    j j �M��`���EP�MQ�M��:&���E������E�M�d�    Y��]� �����������������������������������������U��j�h��d�    P�����3�P�E�d�    �M�M��I��P�M��v���E�    j j �M��f_���E������E�M�d�    Y��]����������������������������U����M��E�P�M�H%��P�M��a��j j �M��^;���MQ�.����P�M���6���E���]� ������������������������U��j�h��d�    P�����3�P�E�d�    �M�E�P�M�Q�M��$�����ra��P�M������E�    j j �M���:���ĊRj �EP�M��'���E������E�M�d�    Y��]� �������������������������������������U��j�h�d�    P�����3�P�E�d�    �M�M���M��P�M��6���E�    j j �M��,:���EP�MQ�M���2���E������E�M�d�    Y��]� ����������������������������������������U��j�hH�d�    P�����3�P�E�d�    �M�M��+M��P�M�����E�    j j �M��9���EP�M��a���E������E�M�d�    Y��]� �����������������������������U��j�hx�d�    P�����3�P�E�d�    �M�M��L��P�M�����E�    j j �M���8���EP�MQ�M���O���E������E�M�d�    Y��]� �����������������������������������������U��j�h��d�    P�����3�P�E�d�    �M�M���K��P�M��f���E�    j j �M��\8���E������E�M�d�    Y��]����������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��-���E�    �M�����UR�M���N���E������E��M�d�    Y��]� ���������������������������������������U��j�h�d�    PQ���3�P�E�d�    �M��EP�M��/-���E�    �M��ȉ�UR�M��5e���E������E��M�d�    Y��]� ���������������������������������������U��j�h8�d�    PQ���3�P�E�d�    �M��EP�M��L4���E�    �M��(��UR�M��c���E������E��M�d�    Y��]� ���������������������������������������U��j�hh�d�    PQ���3�P�E�d�    �M��EP�M��3���E�    �M����UR�M��aY���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��B@���E�    �M��|��UR�M�� 4���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��?���E�    �M��0��UR�M��R���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M���Z���E�    �M��L��UR�M��$���E������E��M�d�    Y��]� ���������������������������������������U��j�h(�d�    PQ���3�P�E�d�    �M��EP�M��XZ���E�    �M��(��UR�M���.���E������E��M�d�    Y��]� ���������������������������������������U��j�hX�d�    PQ���3�P�E�d�    �M��EP�M���0���E�    �M��p��UR�M��q���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��\0���E�    �M��L��UR�M��w���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M���/���E�    �M�����UR�M��#���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��</���E�    �M��h��UR�M��X���E������E��M�d�    Y��]� ���������������������������������������U��Q�M��EPj�MQ�UR�M��B*���E�� ,��E���]� ����������������U��Q�M��EPj �MQ�UR�M��*���E�� ��E���]� ����������������U��Q�M��EPj�MQ�UR�M��:9���E�� ��E���]� ����������������U��Q�M��EPj �MQ�UR�M���8���E�� Č�E���]� ����������������U��j�h�d�    PQ���3�P�E�d�    �M��EP�M��-���E�    �M��x��UR�M��[���E������E��M�d�    Y��]� ���������������������������������������U��j�hH�d�    PQ���3�P�E�d�    �M��EP�M��-���E�    �M��T��UR�M��4���E������E��M�d�    Y��]� ���������������������������������������U��j�hx�d�    PQ���3�P�E�d�    �M��EP�M��,���E�    �M�����UR�M��3���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M���+���E�    �M�����UR�M���K���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��l+���E�    �M�����UR�EP�M��L/���E������E��M�d�    Y��]� ����������������������������������U��j�h�d�    PQ���3�P�E�d�    �M��EP�M���*���E�    �M��؋�UR�EP�M��6���E������E��M�d�    Y��]� ����������������������������������U��j�h8�d�    PQ���3�P�E�d�    �M��EP�M�����E�    �M��l��UR�M��M���E������E��M�d�    Y��]� ���������������������������������������U��j�hh�d�    PQ���3�P�E�d�    �M��EP�M��v���E�    �M��D��UR�M��mW���E������E��M�d�    Y��]� ���������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��,)���E�    �M����j �M����78���E��UR�M���'���E������E��M�d�    Y��]� ��������������������������������������U��j�h��d�    PQ���3�P�E�d�    �M��EP�M��(���E�    �M���j �M����7���E��UR�M�����E������E��M�d�    Y��]� ��������������������������������������U��Q�M��E��M��E���]� ��������U��Q�M��EP�M���'���M��̊�E���]� �����������U��Q�M��EP�M��'���M�����E���]� �����������U��Q�M��EP�M��'���M����E���]� �����������U��Q�M��M���%����]��������������U��Q�M��M��%����]��������������U��Q�M��E�� ���M���6���M�������]�������������U��Q�M��E�� ���M��^���M������]�������������U��Q�M��M��J���M��w����]����������������������U��Q�M��M���'���M��6	����]����������������������U��Q�M��M��_N����]��������������U��Q�M��M��:����]��������������U��Q�M��M��;����]��������������U��Q�M��M������]��������������U��Q�M��M������]��������������U��Q�M��M��t����]��������������U��Q�M�j j�M���K���M��\����]������������������U��Q�M�j j�M���'���M�������]������������������U��Q�M��E�� ���M��m*����]���������������������U��Q�M��E�� ȉ�M��=*����]���������������������U��Q�M��E�� (��M��QR��M�����M��S����]����������������������U��Q�M��E�� ��M��QR�M�����M������]����������������������U��Q�M��E�� |��M��y t�U��BP�kM�����M��QR�\M�����M������]������������������������������U��Q�M��E�� 0��M��y t�U��BP�M�����M��QR��L�����M������]������������������������������U��Q�M��E�� L��M��4����]���������������������U��Q�M��E�� (��M��4����]���������������������U��Q�M��E�� p��M�������]���������������������U��Q�M��E�� L��M������]���������������������U��Q�M��E�� ���M��b����]���������������������U��Q�M��E�� h��M��2����]���������������������U��Q�M��E�� ,��M���?����]���������������������U��Q�M��E�� ��M��?����]���������������������U��Q�M��E�� ��M��+����]���������������������U��Q�M��E�� Č�M�������]���������������������U��Q�M��E�� x��M��B����]���������������������U��Q�M��E�� T��M������]���������������������U��Q�M��E�� ���M�������]���������������������U��Q�M��E�� ���M������]���������������������U��Q�M��E�� ���M���%���M��z����]�������������U��Q�M��E�� ؋�M��A���M��J����]�������������U��Q�M��E�� l��M��1D���M���H����]�������������U��Q�M��E�� D��M��_���M���H����]�������������U��Q�M��E�� ���M����lK���M������]����������U��Q�M��E�� ��M����<K���M������]����������U��Q�M��E��Q��H������]��������U��Q�M��M��K����]��������������U��Q�M��M��+����]��������������U��Q�M��E�� ��M������]���������������������U��Q�M��EP�M��2���E���]� ��������������������U��Q�M��EP�M�����E���]� ��������������������U��Q�M��EP�M���2���M��U�B�A�E���]� ������������������������U��Q�M��EP�M���
���M��U�B�A�E���]� ������������������������U����M��E��;Mtv�M�����} th�U�U��E����t�U����U���E����E��M�+M�M�h-  h<pj�U�R�;������M���U��: t�E�P�MQ�U��P�=�����E���]� ����������������������������������������������U����M��E�;E��   j j�M���C��3�t�U�R�M�����P�M��x.���E�P�M�����P�M�Q�M������P�8�����Ѕ�t,���ĉe�P�M�}�����̉e�Q�M�����M��GC����UR�jB����P�M��68���E���]� ���������������������������������������������������U����M��E�;EtZ�M�Q�M����P�U�R�M�����P�8��������t%3�t!j j�M���B���U�R�M�����P�M��s-���EP�M��$���E���]� ��������������������������������������������U����M��E�;E��   j j�M����3�t�U�R�M�l��P�M�����E�P�M�W��P�M�Q�M��J��P�`-�����Ѕ�t,���ĉe�P�M�k�����̉e�Q�M�@���M��J-����UR�	�����P�M�����E���]� ���������������������������������������������������U����M��E�;EtZ�M�Q�M���P�U�R�M����P�,��������t%3�t!j j�M�����U�R�M�g��P�M�����EP�M��I$���E���]� ��������������������������������������������U����M��E��x t4�MQ�U��J�~��f�E���0��f�E��E�P�M�Q�B������Ѕ�t�E�� �E���]� ���������������������������U����M��E��x t4�MQ�U��J�`��f�E��GF��f�E��E�P�M�Q��@�����Ѕ�t�E�� �E���]� ���������������������������U��Q�M��E��M���E�     �E���]� �������������U����M��EP�M���5���M��U�A;Bu	�E�   ��E�    �E���]� ��������������������U����M��EP�M���%���M��U�A;Bu	�E�   ��E�    �E���]� ��������������������U����M��EP�M��"���ȅ�u	�E�   ��E�    �E���]� ���������������������������U����M��EP�M��9G���ȅ�u	�E�   ��E�    �E���]� ���������������������������U��Q�M��E��H;Msh�  hXohd�������M��K���U�P��]� �������������������U��Q�M��E��H;Msh�  hXohd��������M���	���U�P��]� �������������������U��Q�M��E��H;Msh�  hXohd��{�����M��z+���U�P��]� �������������������U��Q�M��E��H;Msh�  hXohd��+�����M���*���U�P��]� �������������������U��QV�M��M��9����tG�E��x t>�M��$��������M�9Ar'�M�������������M������P�V�M�;Aw_jOhXoh \������ Y��t3�u#hPYh�Yj jPhXoj��������u�j jPhXoh��h�Z�E9�����U��B^��]������������������������������������������������������������U��QV�M��M��9����tG�E��x t>�M��$������)���M�9Ar'�M��������)�����M������P�V�M�;Aw_jOhXoh \������ Y��t3�u#hPYh�Yj jPhXoj��������u�j jPhXohP�h�Z�E8�����U��B^��]������������������������������������������������������������U��Q�M��M������]��������������U��Q�M��M��~6����]��������������U��Q�M��E��H��u�M�������U��: uh�  hЄh8��
�����E�f�@��]�����������������������������U��Q�M��E��H��u�M��C;���U��: uh�  hЄh8��+
�����E�f�@��]�����������������������������U��Q�M��E���]�������������������U��Q�M��E���]�������������������U��QV�M��M�������t0�E��x t'�M���������
�����M������H�N�E�;Pw_jmhXohH��l	����� Y��t3�u#hPYh�Yj jnhXoj�m�������u�j jnhXoh��h�Z�6�����M��Q���E��P�E�^��]�������������������������������������������������������U��QV�M��M��	����t0�E��x t'�M��������&�����M������H�N�E�;Pw_jmhXohH��|����� Y��t3�u#hPYh�Yj jnhXoj�}�������u�j jnhXoh��h�Z�,5�����M��Q���E��P�E�^��]�������������������������������������������������������U��Q�M��E��8 uh  hЄh��������M��+���E���]����������������������������U��Q�M��E��8 uh  hЄh���n�����M������E���]����������������������������U��Q�M��E���]� ����������������U��Q�M��E���]�������������������U��Q�M��E���]� ����������������U��Q�M��E���]�������������������U��Q�M��EP�M��
-���M��U�A+B����]� ���������U��Q�M��EP�M��+���M��U�A+B����]� ���������U��j�h�d�    P�����3�P�E�d�    �M��E�    �E�P�M��c���E�    �MQ�M��9!��P�M�G���U����U��E������M�������E�M�d�    Y��]� ���������������������������������������������U��j�hH�d�    P�����3�P�E�d�    �M��EP�M�Q�M��k@���E�U�U��E�    �M��W7���E��E������M������E�M�d�    Y��]� ������������������������������������������U��j�hx�d�    P�����3�P�E�d�    �M��E�    �E�P�M��i&���E�    �MQ�M������P�M�M&���U����U��E������M�� ���E�M�d�    Y��]� ���������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M��EP�M�Q�M��5����E�U�U��E�    �M��0���E��E������M�������E�M�d�    Y��]� ������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M��E�    �E�P�M������E�    �MQ�M��2��P�M����U����U��E������M��P����E�M�d�    Y��]� ���������������������������������������������U��j�h�d�    P�����3�P�E�d�    �M��E�    �E�P�M��i$���E�    �MQ�M����P�M�M$���U����U��E������M������E�M�d�    Y��]� ���������������������������������������������U��QV�M��M�������tW�E��x tN�M��Q�E�4B�M��x������d��;�r/�M��e������Q�����M��T����H�N�E��H�E�A;�shh�   hXohH�������� Y��t3�u&hPYh�Yj h�   hXoj���������u�j h�   hXoh��h�Z�.�����U��B�M�H�E��P�E�^��]� �����������������������������������������������������������������U��QV�M��M��i�����tW�E��x tN�M��Q�E�4B�M��H��������;�r/�M��5������������M��$����H�N�E��H�E�A;�shh�   hXohH�� ����� Y��t3�u&hPYh�Yj h�   hXoj��������u�j h�   hXoh��h�Z�\-�����U��B�M�H�E��P�E�^��]� �����������������������������������������������������������������U��Q�M��EP�M��\����E���]� ��������������������U��Q�M��EP�M��17���E���]� ��������������������U��Q�M��EP�M��7�����]� �������U��Q�M��EPj�M��9����]� ��������������������U��Q�M��EP�M�������]� �������U��Q�M��EPj�M��������]� ��������������������U��Q�M��E��P�M������]� ���������������������U��Q�M��E��P�M������]� ���������������������U��Q�M��M��3&���E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q��������E���]� ��������������������U��Q�M��M��"���E��t�M�Q�������E���]� ��������������������U��Q�M��M�������E��t�M�Q�A������E���]� ��������������������U��Q�M��M��8���E��t�M�Q�������E���]� ��������������������U��Q�M��M��("���E��t�M�Q��������E���]� ��������������������U��Q�M��M�������E��t�M�Q�������E���]� ��������������������U��Q�M��M��]����E��t�M�Q�A������E���]� ��������������������U��Q�M��M������E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q��������E���]� ��������������������U��Q�M��M��h���E��t�M�Q�������E���]� ��������������������U��Q�M��M��68���E��t�M�Q�A������E���]� ��������������������U��Q�M��M������E��t�M�Q�������E���]� ��������������������U��Q�M��M���"���E��t�M�Q��������E���]� ��������������������U��Q�M��M������E��t�M�Q�������E���]� ��������������������U��Q�M��M�����E��t�M�Q�A������E���]� ��������������������U��Q�M��M��r8���E��t�M�Q�������E���]� ��������������������U��Q�M��M�����E��t�M�Q��������E���]� ��������������������U��Q�M��M�����E��t�M�Q�������E���]� ��������������������U��Q�M��M��X
���E��t�M�Q�A������E���]� ��������������������U��Q�M��M�����E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q��������E���]� ��������������������U��Q�M��M�������E��t�M�Q�������E���]� ��������������������U��Q�M��M�����E��t�M�Q�A������E���]� ��������������������U��Q�M��M��1���E��t�M�Q�������E���]� ��������������������U��Q�M��M�������E��t�M�Q��������E���]� ��������������������U��Q�M��M�����E��t�M�Q�������E���]� ��������������������U��Q�M��M�����E��t�M�Q�A������E���]� ��������������������U��Q�M��M������E��t�M�Q�������E���]� ��������������������U��Q�M��M��3����E��t�M�Q��������E���]� ��������������������U��Q�M��M��)���E��t�M�Q�������E���]� ��������������������U����M��M��Y���j�M��Z���M���M����P�U��P�M��_���M���E����]����������������������������U����M��M������j�M������M���M��-��P�U��P�M������M���E����]����������������������������U����M��E�xs"�M�Q��R�E��P�M���Q�
�����+�U��R�E���P�M�Q�M��]����������U�B    �E��M�Q�P�E��M�Q�Pj j �M��%����]� ���������������������������������������U����M��E�xs"�M�Q��R�E��P�M���Q�O������+�U��R�E���P�M�Q�M������������U�B    �E��M�Q�P�E��M�Q�Pj j �M�����]� ���������������������������������������U����M��E��8 t
�M���U��	�E����E��E���]����������������������U��Q�M���]� ���U��Q�M���]� ���U��Q�M��}u�EP�M������M�HR�u������ �EP�MQ�M��a����U�PP�q������]� ��������������������������������U��Q�M��}u�EP�M������M�HR������ �EP�MQ�M������U�PP�,�������]� ��������������������������������U��QV�M��M�������t�M��������M����;�thh�   hXoh���C���������t3�u&h�h�Yj h�   hXoj�A�������u�j h�   hXoh��hx�������^��]� ���������������������������������������U��QV�M��M��������t�M���������M�����;�thh�   hXoh������������t3�u&h�h�Yj h�   hXoj��������u�j h�   hXoh��hx��-����^��]� ���������������������������������������U��j�h0�d�    PQ�� SVW���3�P�E�d�    �e��M�E���E�M����;E�s�M�M��R�E�3ҹ   ��U�J��;�w�8�U�r��M��Q��+ƋM�9Aw�U�B��M�A�E���M��,���E��E�    �U�R�M�������E܋E��P�M������E؋M؉M��g�e��U�U��E��E�P�M������EԋM��Q�M��j����EЋUЉU��j j�M��Q!��j j �%����F��E�   ��E�   ��F��E�������E������} v�EP�M������P�M�Q������j j�M��� ���U�R�E��P�M�Q�M��������m���U�E�B�MQ�M��p���M�d�    Y_^[��]� ������������������������������������������������������������������������������������������������������������������������U��j�h`�d�    PQ�� SVW���3�P�E�d�    �e��M�E���E�M��g���;E�s�M�M��R�E�3ҹ   ��U�J��;�w�8�U�r��M��0���+ƋM�9Aw�U�B��M�A�E���M������E��E�    �U�R�M������E܋E��P�M������E؋M؉M��g�e��U�U��E��E�P�M��u����EԋM��Q�M�������EЋUЉU��j j�M��w���j j ������H��E�   ��E�   ��H��E�������E������} v�EP�M����P�M�Q�������j j�M������U�R�E��P�M�Q�M�������������U�E�B�MQ�M�������M�d�    Y_^[��]� ������������������������������������������������������������������������������������������������������������������������U������3ŉE��M��E�    �E��P�M�Q�UR�E�P�)������t�M�M���   k� �L�M�E�M�3��:�����]� ���������������������������U������3ŉE��M��E�    �E��P�M�Q�UR�E�P�*)������t�M�M���   k� �L�M�E�M�3�������]� ���������������������������U����M��E�    �E��P�M�Qj�UR�E�P�(������}���  f�M��f�U�f�U�f�E���]� ����������������������������������U����M��E�    �E��P�M�Qj�UR�E�P�(������}���  f�M��f�U�f�U�f�E���]� ����������������������������������U����M��E��8 u	�E�   ��E�    �E���]�������������������������U����M�3�f�E��M��U�Q�E�P�M������M�HR��������]� �����������������������U����M�3�f�E��M��U�Q�E�P�M��	���M�HR���������]� �����������������������U����E�E�M��%�U���U�E�� t�M��+�U���U�E��t�M��#�U���U�E�� .�M���M�U��*�E���E��M��t�U�E��M���M�U�� 0  �U��E��tP�}�    u�E�f�.�}� 0  u�E�A��}�   u�E�E��E�G�M��M��U��U��E�M���U���U��N�}�    u�E�f�.�}� 0  u�E�a��}�   u�E�e��E�g�E��E��M��M��U�E���M���M�U�� �E��]����������������������������������������������������������������������������������U����E�E�M��%�U���U�E�� t�M��+�U���U�E��t�M��#�U���U�E�� .�M���M�U��*�E���E��M��t�U�E��M���M�U�� 0  �U��E��tP�}�    u�E�f�.�}� 0  u�E�A��}�   u�E�E��E�G�M��M��U��U��E�M���U���U��N�}�    u�E�f�.�}� 0  u�E�a��}�   u�E�e��E�g�E��E��M��M��U�E���M���M�U�� �E��]����������������������������������������������������������������������������������U��j�h��d�    P���   ���3ŉE�VP�E�d�    h`  h���EP�������}0 v�M ���+t�E ���-u	�E�   ��E�    �U��U��M�q��% 0  = 0  tǅ|���X��Jǅ|���\��E���;E0w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M���|���R�   k� M Q�������E�f�`�f�U�������   k� � �   k� ��T��   k� �T�R�   k� M Q�u�����E���`���R�M�*�����l�����l�����\����E�    ��\���Q������E��E�������`��������j0�M������f�E�j �U0R�M�������E�   j �M�����P�E E0P�   k� U R�M������p���P�M������d�����d�����h����E���h���R��������E��E���p����N����E�P�M�������E��M��j
��f�E��M$�M��U�;U0u �E�E��E��M�Q�U$R�E�P�M��W���e�M�M��M��U�R�E,P�M�Q�M��7���U�R�E(P�M���Q�M�����M����f���U�R�M�����f�0�E�P�M$Q�U�R�M�����j �M������E��E����tY�U����~O�M���E�+E�;�s?�M���E�+E��M�Qj�U�R�M�����   �� �M����~	�E����E�뜍M��K���E0�M�������t�����x�����x��� |(	��t��� v�M�����;E0v�M����+E0�E���E�    �M��M��M�D��%�  �E��}�@ty�}�   tp�U�R�EP�MQ�UR��<���P�MQ�<������@�U�E�E�    �M�Qj �M��W���P�UR�EP��T���Q�UR���������P�M�U�   �}�   um�E�Pj �M�����P�MQ�UR��,���P�MQ��������@�U�E�M�Q�UR�EP�MQ��D���R�EP�������P�M�U�E�    �5�E�Pj �M�����P�MQ�UR��4���P�MQ�1�������@�U�E�M0+M�Q�U�R�M��m���P�EP�MQ��L���R�EP���������P�M�Uj j �M�����E�P�MQ�UR�EP�MQ�UR�������E��M������E������M������E�M�d�    Y^�M�3��C�����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h&�d�    P���   ���3ŉE�VP�E�d�    h`  h���EP�4�����}0 v�M ���+t�E ���-u	�E�   ��E�    �U��U��M���% 0  = 0  tǅ|���X��Jǅ|���\��E���;E0w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M���|���R�   k� M Q�������E�f�`�f�U�������   k� � �   k� ��T��   k� �T�R�   k� M Q������E���`���R�M�J�����l�����l�����\����E�    ��\���Q�������E��E�������`��������j0�M����f�E�j �U0R�M�����E�   j �M��?���P�E E0P�   k� U R�M�������p���P�M������d�����d�����h����E���h���R�
������E��E���p����n����E�P�M��7����E��M��k���f�E��M$�M��U�;U0u �E�E��E��M�Q�U$R�E�P�M������e�M�M��M��U�R�E,P�M�Q�M��j����U�R�E(P�M���Q�M��R����M�����f���U�R�M��F���f�0�E�P�M$Q�U�R�M��#���j �M��:����E��E����tY�U����~O�M���E�+E�;�s?�M���E�+E��M�Qj�U�R�M�������   �� �M����~	�E����E�뜍M�����E0�M������t�����x�����x��� |(	��t��� v�M�����;E0v�M�����+E0�E���E�    �M��M��M�d��%�  �E��}�@ty�}�   tp�U�R�EP�MQ�UR��<���P�MQ��������@�U�E�E�    �M�Qj �M������P�UR�EP��T���Q�UR��������P�M�U�   �}�   um�E�Pj �M�����P�MQ�UR��,���P�MQ���������@�U�E�M�Q�UR�EP�MQ��D���R�EP�������P�M�U�E�    �5�E�Pj �M��M���P�MQ�UR��4���P�MQ�l�������@�U�E�M0+M�Q�U�R�M�����P�EP�MQ��L���R�EP�2�������P�M�Uj j �M�!����E�P�MQ�UR�EP�MQ�UR�c�����E��M������E������M��G����E�M�d�    Y^�M�3��c�����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��M��y����M������E��Q�M������j�U��P�M�����M��    ��]�����������������������������U����M��M������M��<����E��Q�M�����j�U��P�M�����M��    ��]�����������������������������U��Q�M��M����E��]� ��������U��Q�M��M������E��]� ��������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �8����E�h^  h��M�Qj4�������E��E�    �}� t:j �M����P�M������E��U��U��E��E����E��M�Q�M���	���E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�hs  h��M�Qj4�_������E��E�    �}� t:j �M�����P�M��u����E��U��U��E��E����E��M�Q�M�����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��x���3ŉE�P�E�d�    �E�    �} ��   �E�8 ��   �����E�jChX��M�Qj�������E��E�    �}� tbj �U�R�M�s����E��E��E��E��MЃ��MЋM������P��|��������E��U��U��E�   �EЃ��EЋM�Q�M������E���E�    �UȉU��E�   �E�M���E�   �UЃ�t�e����|����"���E������EЃ�t�e���M������   �M�d�    Y�M�3��6�����]������������������������������������������������������������������������������������������U��j�h-�d�    P��x���3ŉE�P�E�d�    �E�    �} ��   �E�8 ��   �����E�jChX��M�Qj�������E��E�    �}� tbj �U�R�M������E��E��E��E��MЃ��MЋM��\���P��|����p����E��U��U��E�   �EЃ��EЋM�Q�M�����E���E�    �UȉU��E�   �E�M���E�   �UЃ�t�e����|�������E������EЃ�t�e���M�������   �M�d�    Y�M�3�������]������������������������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �x����E�hO  h��M�QjD��������E��E�    �}� t:j �M�_���P�M�������E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��
���   �M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �8����E�hl
  h��M�QjD�������E��E�    �}� t:j �M����P�M������E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�jMh��M�Qj�b������E��E�    �}� t:j �M�����P�M��x����E��U��U��E��E����E��M�Q�M��\����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]�����������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�jMh��M�Qj�"������E��E�    �}� t:j �M����P�M��8����E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��P���   �M�d�    Y��]�����������������������������������������������������������������������������U��j�hD�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �x����E�h�  h��M�Qj��������E��E�    �}� t:j �M�_���P�M�������E��U��U��E��E����E��M�Q�M��M����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �8����E�h�  h��M�Qj�������E��E�    �}� t:j �M����P�M������E��U��U��E��E����E��M�Q�M��Y����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h$�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�h�  h��M�Qj�_������E��E�    �}� t:j �M�����P�M��u����E��U��U��E��E����E��M�Q�M��D����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h�  h��M�Qj�������E��E�    �}� t:j �M����P�M��5����E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��M���   �M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �x����E�h(  h��M�QjX��������E��E�    �}� t<jj �M�]���P�M�������E��U��U��E��E����E��M�Q�M��!����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�� ���   �M�d�    Y��]������������������������������������������������������������������������U��j�ht�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �8����E�h(  h��M�QjX�������E��E�    �}� t<jj �M����P�M������E��U��U��E��E����E��M�Q�M�����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�������   �M�d�    Y��]������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�h(  h��M�QjX�_������E��E�    �}� t<jj �M�����P�M��s����E��U��U��E��E����E��M�Q�M��L����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]������������������������������������������������������������������������U��j�hT�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h(  h��M�QjX�������E��E�    �}� t<jj �M����P�M��3����E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��K����   �M�d�    Y��]������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �x����E�h  h���M�Qj��������E��E�    �}� t:j �M�_���P�M�������E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h4�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �8����E�h  h���M�Qj�������E��E�    �}� t:j �M����P�M������E��U��U��E��E����E��M�Q�M�萾���E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�hD  h���M�Qj�_������E��E�    �}� t:j �M�����P�M��u����E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�hD  h���M�Qj�������E��E�    �}� t:j �M����P�M��5����E��U��U��E��E����E��M�Q�M��	����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��M����   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �x����E�h�   h���M�Qj�߼�����E��E�    �}� t<jj �M�]���P�M�������E��U��U��E��E����E��M�Q�M��-����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �8����E�h�   h���M�Qj蟻�����E��E�    �}� t<jj �M����P�M������E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�������   �M�d�    Y��]������������������������������������������������������������������������U��j�hd�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�h�   h���M�QjD�_������E��E�    �}� t:j �M�����P�M��u����E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h�   h���M�QjD�������E��E�    �}� t:j �M����P�M��5����E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��M����   �M�d�    Y��]��������������������������������������������������������������������������U��j�hD�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �x����E�h  h���M�Qj�߷�����E��E�    �}� t:j �M�_���P�M�������E��U��U��E��E����E��M�Q�M��=����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h��d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �8����E�h|  h���M�Qj蟶�����E��E�    �}� t:j �M����P�M������E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�������   �M�d�    Y��]��������������������������������������������������������������������������U����M��}����E�U��E�M��U��P�E��]� ���������������������U��Q�M�������]�����������������U����M��5����E��}� t�E�P�M��������M�Q�������M��������Ѕ�u�M����?����E���E����E��]�������������������������������U��j�h�d�    P��   ���3ŉE�VP�E�d�    �M�����% 0  = 0  u%�EP�MQ�UR�EP�MQ�UR�g�������  ��L���P�M�.�����\�����\�����T����E�    ��T���R�l�������p����E�������L����ޠ���E�P��p����~����E�   �M�M��E� ��P���R�M������X�����X�����`����E���`���Q��������h����E���P����u����U�R�   k�����Q�   k� ��P��h����p����MQ�UR�����������t�h�M脼���Ⱥ   k��T�;�u�E�� +�M����M��M������3�M�O����и   k�
�D�;�u�M��-�U����U��M�����E� �E�    �E�    j �M��1�����|�����|������t��|��������   ��E��M�m����MQ�UR�����������te�M趻����Q�U�R�������E��}�
sD�}�$|�E����E��.�}� u�}� u� �M��U�������M����M��U����U��x����;  �M��D�����u3�f��v������p����
���f��v���f��v���f��x���j j�M��´���E��E�    ��M�����UR�EP�������ȅ���   �M�ٺ����R�E�P�������E��}�
s~�E��}�$|�M����M��.�}� u�}� u� �U��E������
�U����U��E����E��M�Q�M��7������t%�E�P�M��#�����l�����l��������l�����M�M�Q�M���������t!��x�����t�M��������x���;�t��j j�M������E����E�������}� u�"�M�Q�M�袨�����~�E����E���E��M�����   �}� ��   ��|������u�{�t�M����M�t��|����2�E�P�M��D����;�u"�}� u"��|����2�E�P�M��"����;�}�E��%�   �� ��|������~��|�������|����_����E��M��8����E���t�}� u�M��0�U����U��EP�MQ�������Ѕ�tE�M�ݸ������p���������;�u(�׳���   k� � �M����E����E��M�8����}� uj��E��M�$����MQ�UR����������t'�M�m����Ⱥ   k� �T�;�u�E����E�붃}� }�M��0�U����U��E����E���E��M�����MQ�UR�:���������tI�M������Q�U�R��������E��}�
s(�}�$} �E��M�������E����E��M����M���U�����  �EP�MQ��������Ѕ���  �M蓷�����   k��L�;�t �M�w����и   k��D�;��i  �M��e�U����U��M������E� �E�    �EP�MQ�������Ѕ�t�h�M�������   k��L�;�u�U��+�E����E��M�����3�M�����Ⱥ   k�
�T�;�u�E�� -�M����M��M�T����UR�EP��������ȅ�t*�M蝶���и   k� �D�;�u�E��M������M���t�U��0�E����E���E��M������MQ�UR�n���������tI�M�7�����Q�U�R�������E��}�
s(�}�} �E��M�������E����E��M����M���U���u�E���u�M�M��U�� �E���d����E������M�������d����M�d�    Y^�M�3�葻����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��   ���3ŉE�VP�E�d�    �M�y���% 0  = 0  u%�EP�MQ�UR�EP�MQ�UR��������  ��L���P�M�ν����\�����\�����T����E�    ��T���R� �������p����E�������L����~����E�P��p����D����E�   �M�M��E� ��P���R�M�_�����X�����X�����`����E���`���Q跘������h����E���P��������U�R�   k����Q�   k� �P��h��������MQ�UR蟠��������t�h�M�3����Ⱥ   k��T�;�u�E�� +�M����M��M������3�M������и   k�
�D�;�u�M��-�U����U��M�����E� �E�    �E�    j �M��ѡ����|�����|������t��|��������   ��E��M�L����MQ�UR�X���������te�M�e�����Q�U�R�\������E��}�
sD�}�$|�E����E��.�}� u�}� u� �M��U������M����M��U����U��x����;  �M�������u3�f��v������p���苘��f��v���f��v���f��x���j j�M��b����E��E�    ��M�s����UR�EP�������ȅ���   �M������R�E�P�������E��}�
s~�E��}�$|�M����M��.�}� u�}� u� �U��E�����
�U����U��E����E��M�Q�M��מ�����t%�E�P�M��Þ����l�����l��������l�����M�M�Q�M�蜞�����t!��x�����t�M���������x���;�t��j j�M�躬���E����E�������}� u�"�M�Q�M��B������~�E����E���E��M�����   �}� ��   ��|������u�{�t�M����M�t��|����2�E�P�M������;�u"�}� u"��|����2�E�P�M�����;�}�E��%�   �� ��|������~��|�������|����_����E��M��أ���E���t�}� u�M��0�U����U��EP�MQ�������Ѕ�tE�M��������p���������;�u(�w����   k� � �M����E����E��M�����}� uj��E��M�����MQ�UR����������t'�M�����Ⱥ   k� �T�;�u�E����E�붃}� }�M��0�U����U��E����E���E��M�����MQ�UR襮��������tI�M������Q�U�R�������E��}�
s(�}�$} �E��M������E����E��M����M���U�����  �EP�MQ�9������Ѕ���  �M�B������   k��L�;�t �M�&����и   k��D�;��i  �M��e�U����U��M�����E� �E�    �EP�MQ�7������Ѕ�t�h�M��������   k��L�;�u�U��+�E����E��M�h����3�M�����Ⱥ   k�
�T�;�u�E�� -�M����M��M�3����UR�EP�?������ȅ�t*�M�L����и   k� �D�;�u�E��M�������M���t�U��0�E����E���E��M������MQ�UR�٬��������tI�M������Q�U�R��������E��}�
s(�}�} �E��M������E����E��M����M���U���u�E���u�M�M��U�� �E���d����E������M�聠����d����M�d�    Y^�M�3��1�����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P���   ���3ŉE�VP�E�d�    ��0���P�M觳����@�����@�����8����E�    ��8���R��������T����E�������0����W����E�P��T���������E�   ��4���Q�M�B�����<�����<�����D����E���D���P�7�������L����E���4���������M�Q�   k�(�P�   k� ��(�R��L���������E��x���ƅw��� �MQ�UR�i���������t�z�M������Ⱥ   k��T�;�u"��x���� +��x�������x����M�[����<�M蹧���и   k��D�;�u ��x����-��x�������x����M������x���� 0��x�������x�����x����x��x�������x���ƅ��� ǅp���    ǅd���    �MQ�UR苲��������u�M�����Ⱥ   k� �T�;�t�e�EP�M葹��P�������ȅ�tB�M�����и   k��D�;�t�M�Ŧ���Ⱥ   k��T�;�u
�M�A����ƅ���j �M�迖����`�����`������t��`��������   �ƅ����M������MQ�UR�x�����������   �M�=�����Q�U�R��������h�����h���se��p���$|��d�������d����F��h��� u��p��� u�2��x�����h�����(����x�������x�����p�������p����J����  �M�褞����u3�f��Z������T����j���f��Z���f��Z���f��\���j j�M��"����E�ǅl���    ��M�����UR�EP�q������ȅ��.  �M�6�����R�E�P��������h�����h�����   ƅ�����p���$|��d�������d����F��h��� u��p��� u�2��x�����h�����(��
��x�������x�����p�������p�����l���Q�M��c������t(��l���P�M��L�����P�����P��������P�����V��l���Q�M��"������t!��\�����t�M�B�������\���;�t�"�j j�M��@�����l�������l���������l��� u�.��l���Q�M�輒�����~��l�������l����ƅw�����w�������   ��l��� ��   ��`������u
�   �   ��l�������l���t��`����2��l���P�M��@����;�u(��l��� u(��`����2��l���P�M������;�}	ƅw����%�   �� ��`������~��`�������`����A����E��M��+����������t!��p��� u��x����0��x�������x����EP�MQ��������Ѕ�tN�M���������T���������;�u1軝���   k� � ��x�������x�������x����M������p��� ��   �ƅ����M������MQ�UR�u���������t-�M�>����Ⱥ   k� �T�;�u��d�������d���뭃�d��� }'��x����0��x�������x�����d�������d����ƅ����M�p����MQ�UR�����������tg�M蹡����Q�U�R��������h�����h���s@��p���$}2��x�����h�����(����x�������x�����p�������p����s�����������  �EP�MQ�c������Ѕ���  �M�(������   k��L�;�t �M�����и   k��D�;���  ��x����p��x�������x����M�l���ƅ��� ǅp���    �EP�MQ�������Ѕ�t�z�M袠�����   k��L�;�u"��x����+��x�������x����M�����<�M�d����Ⱥ   k��T�;�u ��x���� -��x�������x����M�Ȳ���UR�EP�H������ȅ�t-�M�����и   k� �D�;�uƅ����M膲����������t��x����0��x�������x����ƅ����M�P����MQ�UR�����������tg�M號����Q�U�R�w�������h�����h���s@��p���}2��x�����h�����(����x�������x�����p�������p����s�����w�����u�������u	�M��x�����x���� �E��d����ǅH���    �E������M�������H����M�d�    Y^�M�3�轤����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hf�d�    P���   ���3ŉE�VP�E�d�    ��0���P�M触����@�����@�����8����E�    ��8���R��������T����E�������0����W���E�P��T��������E�   ��4���Q�M�B�����<�����<�����D����E���D���P蚁������L����E���4�����~���M�Q�   k�ܒP�   k� ��ܒR��L����ǒ���E��x���ƅw��� �MQ�UR�r���������t�z�M�����Ⱥ   k��T�;�u"��x���� +��x�������x����M�����<�M�Ȯ���и   k��D�;�u ��x����-��x�������x����M�\�����x���� 0��x�������x�����x����x��x�������x���ƅ��� ǅp���    ǅd���    �MQ�UR蔈��������u�M�*����Ⱥ   k� �T�;�t�e�EP�M�����P�������ȅ�tB�M�����и   k��D�;�t�M�ԭ���Ⱥ   k��T�;�u
�M�����ƅ���j �M�迉����`�����`������t��`��������   �ƅ����M�7����MQ�UR�C�����������   �M�L�����Q�U�R�C�������h�����h���se��p���$|��d�������d����F��h��� u��p��� u�2��x�����h�����ܒ���x�������x�����p�������p����J����  �M�褑����u3�f��Z������T����K���f��Z���f��Z���f��\���j j�M��"����E�ǅl���    ��M�0����UR�EP�<������ȅ��.  �M�E�����R�E�P�<�������h�����h�����   ƅ�����p���$|��d�������d����F��h��� u��p��� u�2��x�����h�����ܒ�
��x�������x�����p�������p�����l���Q�M��c������t(��l���P�M��L�����P�����P��������P�����V��l���Q�M��"������t!��\�����t�M�Q�������\���;�t�"�j j�M��@�����l�������l���������l��� u�.��l���Q�M�輅�����~��l�������l����ƅw�����w�������   ��l��� ��   ��`������u
�   �   ��l�������l���t��`����2��l���P�M��@����;�u(��l��� u(��`����2��l���P�M������;�}	ƅw����%�   �� ��`������~��`�������`����A����E��M��+����������t!��p��� u��x����0��x�������x����EP�MQ�Ö�����Ѕ�tN�M�Щ������T����������;�u1軐���   k� � ��x�������x�������x����M�R�����p��� ��   �ƅ����M�4����MQ�UR�@���������t-�M�M����Ⱥ   k� �T�;�u��d�������d���뭃�d��� }'��x����0��x�������x�����d�������d����ƅ����M诽���MQ�UR軕��������tg�M�Ȩ����Q�U�R迳������h�����h���s@��p���$}2��x�����h�����ܒ���x�������x�����p�������p����s�����������  �EP�MQ�.������Ѕ���  �M�7������   k��L�;�t �M�����и   k��D�;���  ��x����p��x�������x����M諼��ƅ��� ǅp���    �EP�MQ�������Ѕ�t�z�M豧�����   k��L�;�u"��x����+��x�������x����M�E����<�M�s����Ⱥ   k��T�;�u ��x���� -��x�������x����M�����UR�EP�������ȅ�t-�M� ����и   k� �D�;�uƅ����M�Ż����������t��x����0��x�������x����ƅ����M菻���MQ�UR蛓��������tg�M訦����Q�U�R蟱������h�����h���s@��p���}2��x�����h�����ܒ���x�������x�����p�������p����s�����w�����u�������u	�M��x�����x���� �E��d����ǅH���    �E������M�������H����M�d�    Y^�M�3�轗����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M��E�P�M讙���E�M�M��E�    �U�R謥�����E��E������M��pr���	�E(���E(�M(�����   �E(���%uO�U(���U(j �E(�Q�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M���M��B$�Ћ�P�M�U�   �E(��� uB��M�ܠ���UR�EP�\������ȅ�t�M�%�����RjH�M�萺������t���<j �M������Q�M�螐���ЋE(�;�t�U ����M ����M�h��������UR�EP�������ȅ�t�U ����M ��U�E��M�J�E�M�d�    Y��]�$ �����������������������������������������������������������������������������������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M��E�P�M莗���E�M�M��E�    �U�R��r�����E��E������M��Pp���	�E(���E(�M(�����   �E(���%uO�U(���U(j �E(�Q�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M���M��B$�Ћ�P�M�U�   �E(��� uB��M������UR�EP�������ȅ�t�M������RjH�M��-�������t���<j �M������Q�M���t���ЋE(�;�t�U ����M ����M致�������UR�EP�z�����ȅ�t�U ����M ��U�E��M�J�E�M�d�    Y��]�$ �����������������������������������������������������������������������������������������������������������������������U��j�h �d�    P���   ���3ŉE�VP�E�d�    �EP�Л������X����M�Q��X���������E�    �M�芃����u3�f��f������X����P���f��f���f��f���f��h����MQ�%�������8����U�R�   k�����Q�   k� ��P��8��������M��|����UR�EP�m������ȅ�t�z�M������и   k��D�;�u"��|����+��|�������|����M�_����<�M轉�����   k��L�;�u ��|����-��|�������|����M�!����M��   �M�}   uǅ`���   �I�}   uǅD���   �(�} uǅL���    �
ǅL���
   ��L�����D�����D�����`�����`�����p����E� ƅw��� �UR�EP� ������ȅ���   �M�����и   k� �D�;���   �E��M�Y����MQ�UR�ٸ��������tb�M袈���Ⱥ   k��T�;�t�M膈�����   k��L�;�u*��p��� t	��p���uǅp���   �E� �M�������p��� u
ǅp���   ��p��� t6��p���
t-��p���uǅT���   �
ǅT���   ��T�����H����
ǅH���
   ��H�����@����M�Qj�M�肁���E�ǅx���    �   k�E��<�����M�@����MQ�UR������������!  �M腇����Q�U�R�c�������P�����P���;�@�����   ��|�����P����������w�����u��|������0t$��|���;�<���s��|�������|���ƅw����E���x���P�M��u�����t(��x���R�M��u����\�����\��������\����
�V��x���P�M��~u�����t!��h�����t�M螆������h���;�t�"�j j�M�蜃����x�������x���������x��� u�+��x���P�M��u�����~��x�������x�����E� j �M��Uv����l����E�����   ��x��� ��   ��l������u
�   �   ��x�������x���t��l����1��x���R�M��t��� ;�u(��x��� u%��l����1��x���R�M��jt��� ;�}�E� �%�   �� ��l����
��~��l�������l����G����U���t%��w�����u��|����0��|�������|�����E���u	�M��|�����|���� ��p�����4����E� �M��-z���E������M��z����4����M�d�    Y^�M�3��Ί����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hp�d�    P���   ���3ŉE�VP�E�d�    �EP�Dg������X����M�Q��X����z����E�    �M���{����u3�f��f������X����j��f��f���f��f���f��h����MQ��h������8����U�R�   k����Q�   k� �P��8����$z���M��|����UR�EP��p�����ȅ�t�z�M�j����и   k��D�;�u"��|����+��|�������|����M������<�M�,������   k��L�;�u ��|����-��|�������|����M������M��   �M�}   uǅ`���   �I�}   uǅD���   �(�} uǅL���    �
ǅL���
   ��L�����D�����D�����`�����`�����p����E� ƅw��� �UR�EP�K������ȅ���   �M�T����и   k� �D�;���   �E��M������MQ�UR����������tb�M�����Ⱥ   k��T�;�t�M��������   k��L�;�u*��p��� t	��p���uǅp���   �E� �M聩�����p��� u
ǅp���   ��p��� t6��p���
t-��p���uǅT���   �
ǅT���   ��T�����H����
ǅH���
   ��H�����@����M�Qj�M���y���E�ǅx���    �   k�E��<�����M�ߨ���MQ�UR�����������!  �M�������Q�U�R��������P�����P���;�@�����   ��|�����P���������w�����u��|������0t$��|���;�<���s��|�������|���ƅw����E���x���P�M��n�����t(��x���R�M��n����\�����\��������\����
�V��x���P�M���m�����t!��h�����t�M��������h���;�t�"�j j�M���{����x�������x���������x��� u�+��x���P�M��xm�����~��x�������x�����E� j �M��n����l����E�����   ��x��� ��   ��l������u
�   �   ��x�������x���t��l����1��x���R�M���l��� ;�u(��x��� u%��l����1��x���R�M���l��� ;�}�E� �%�   �� ��l����
��~��l�������l����G����U���t%��w�����u��|����0��|�������|�����E���u	�M��|�����|���� ��p�����4����E� �M��r���E������M��~r����4����M�d�    Y^�M�3��.�����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���@���3ŉE��E܉EԋMQ�UR����������t�[j �M�u{����Q�M �~���E��Uۃ�+u�E�� +�Mԃ��MԋM�ލ��� �Uۃ�-u�E�� -�Mԃ��MԋM輍���E� �UR�EP�8������ȅ�t,j �M��z����R�M �}������0u�E��M�w�����Mڅ�t�U��0�Eԃ��EԹ   k��D܉E���E��M�A����MQ�UR�����������tFj �M�z����Q�M �$}���E��Uۃ�0|$�Eۃ�9�MԊUۈ�E�;E�s	�Mԃ��M���Uڅ�u�E܉EԋM�� �E�    �U�Rj
�E�P�M�Q赃�����E��E�    �UR�EP�b������ȅ�t	�UЃ��UЍE�9E�t�}� u�M�;M|�U;U�}�EЃ��E���M�Ủ�EЋM�3������]����������������������������������������������������������������������������������������������������������������������������������U���@���3ŉE��E܉EԋMQ�UR�rg��������t�[j �M������Q�M ��a���E��Uۃ�+u�E�� +�Mԃ��MԋM蝡��� �Uۃ�-u�E�� -�Mԃ��MԋM�{����E� �UR�EP�y�����ȅ�t,j �M莌����R�M �qa������0u�E��M�6�����Mڅ�t�U��0�Eԃ��EԹ   k��D܉E���E��M� ����MQ�UR�y��������tFj �M������Q�M ��`���E��Uۃ�0|$�Eۃ�9�MԊUۈ�E�;E�s	�Mԃ��M���Uڅ�u�E܉EԋM�� �E�    �U�Rj
�E�P�M�Q�5������E��E�    �UR�EP��e�����ȅ�t	�UЃ��UЍE�9E�t�}� u�M�;M|�U;U�}�EЃ��E���M�Ủ�EЋM�3��}����]����������������������������������������������������������������������������������������������������������������������������������U��j�h
�d�    P���  ���3ŉE�VP�E�d�    ��t���ǅ|���    h�  h(��E�HQ�R�E�HQ�R�)������E��tQ������Q�M������������������ ����E�    �� ���P�2|������p����E������������Y���O������Q�M蘀���������������������E�   ������P�?�������p����E������������HY��ƅ���� ƅw��� �M��O����E�   ��4���Q��p����d���M��h����E�������R�M�����������������������E�������Q��������$����E���������X���UR�   k���̒Q�   k� ̒P��$���迚��ǅ`���    ���`�������`������������K  ��`����>  ��`�����4�����<�����<����� ��<�����<���X�	  ��<�����T��$�@��U�R��p����k����E�������BV���E��M�n�����u=�EP�MQ�b������Ѕ�t&�M�+t�����M����� ;�tj �M��y���Q��`���uH�M��ť����w;�MQ�UR�H��������u�M��s�����M��~���;�t
j �M��Hy����h���R�M��k���������������������E�������Q�������s���E���h����g_��������赐���M������UR�EP�y������ȅ�tv��\���R�M��\��������������x����E���|�������|�����x���R������q�������t)�M��r�����������k���;�uǅ(���   �
ǅ(���    ��(�����^����E�   ��|�����t��|������\����^����^�����t������D���R�M���[���������������������E�	������Q������������\����E���D����/^����\�����tƅ�����E�������Y^���E��M��Hh���  �EP�MQ�]}�����Ѕ�t�t  ������P��p����T���������������������E�
��|�������|����������w�����vej ������P��p����TT���������������������E�   ��|�������|�����������k���0�M�Xq����;�uǅ���   �
ǅ���    �������Z����E�
   ��|�����t��|�����������Bg���E�   ��|�����t��|�����������g����Z�����t?�M�l���������R��p����S��������������P�M��i����������f���!  �����Q��p����:����������������������E���|�������|����������$�����vej ������Q��p��������������������������E�   ��|�������|����������j���0�M�p����;�uǅ���   �
ǅ���    �������S����E�   ��|�����t��|���������e���E�   ��|�����t��|�����������e����S�����tF�M������H���P��p������������������Q�M��g����H����e��ƅw�����   ��,���R��p�����Q��������������������uǅ ���   �
ǅ ���    �� �����_�����,����&e����_�����t�f������R��p����~��������������舠����uǅ,���   �
ǅ,���    ��,�����[�����������d����[�����tƅw�����  ǅT���    ��p����Co����8�����d���R��p���赅���E���d����3g����u3�f��B������p����Dx��f��B���f��B���f��H�����H�����t��d����]��� ��|e��M�|����MQ�UR�����������t?�M��m����Q�UR裠������h�����h���
s��h�����̒Q�M���\����M  j j�M��.g���E�ǅx���    ��M�����UR�EP�}������ȅ���   �M�Bm����R�EP� �������h�����h���
sW��h�����̒R�M��U\����x���P�M���[�����t(��x���R�M��[���������������������
�K��x���P�M��[�����t�M�l������H���;�t�"�j j�M��i����x�������x���������x��� u�.��x���R�M��([��� ��~��x�������x����ƅ������d����D[����L�������������   ��x��� ��   ��L������u
�   �   ��x�������x���t��L����0��x���Q�M��Z���;�u(��x��� u(��L����0��x���Q�M��sZ���;�}	ƅ�����%�   �� ��L������~��L�������L����A�����������t �E��M��{`���E���d����l`����  �E��M��[`����p����6���f��D����UR�EP�B������ȅ���   ��D�������   �M��j������D���;���   �UR�M�r}��P�����������t\��T���;�8���}N�M�j����R�EP蒝������h�����h���
s'��h�����̒R�M���Y����T�������T���눋�T���;�8���}ƅ�����M��Ic����u	ƅ�����+���T�������T�����T���;�8���}j0�M��cY�����E���d����)_���   ��`���u�vƅo��� ��M�|���MQ�UR����������t)�M��i����QjH��$����2����Ѕ�t	ƅo���븋�`�����4����� u��o�����uƅ������������������  �M��1�������  �������;K���E���,���Q�M��!a���������������������E�������P�������i���E���,�����T����M�{����P���Q�M��DR����������������|����E���|����� ��|�����|���Q������������� ~���Ѕ�t@�EP�MQ�Ę�����Ѕ�t)�M�h�����������a��� ;�uǅ0���   �
ǅ0���    ��0�����]����E�   ��|����� t��|���ߍ�P����#T����]�����t������8���Q�M��fQ���������������������E�������P�������X}����g����E���8�����S����g�����tƅ�����E���������S����������tj �M��C������w�����tj-jj �M��̘���M�Q�M�/\����|�����@��|����E��M��}\���E������M��]���E�M�d�    Y^�M�3��!m����]� ��i���b�����  �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P���  ���3ŉE�VP�E�d�    ��t���ǅ|���    h�  h(��E�HQ�R�E�HQ�R��~�����E��tQ������Q�M��l���������������� ����E�    �� ���P藋������p����E������������E���O������Q�M�l���������������������E�   ������P�P������p����E������������XE��ƅ���� ƅw��� �M��v���E�   ��4���Q��p���迆���M��x����E�������R�M�l���������������������E�������Q�vG������$����E���������D���UR�   k�����Q�   k� ��P��$����X��ǅ`���    ���`�������`������������K  ��`����>  ��`�����4�����<�����<����� ��<�����<���X�	  ��<�����D��$�0��U�R��p����Zb���E�������a���E��M�~�����u=�EP�MQ�=a�����Ѕ�t&�M�Jt�����M��y{��� ;�tj �M��m����Q��`���uH�M�������w;�MQ�UR�aN��������u�M��s�����M��&{���;�t
j �M�������h���R�M��,����������������������E�������Q������@Z���E���h�����S��������������M�H����UR�EP�T`�����ȅ�tv��\���R�M��S��������������x����E���|�������|�����x���R�������b������t)�M�s���������薃���;�uǅ(���   �
ǅ(���    ��(�����^����E�   ��|�����t��|������\�����R����^�����t������D���R�M��LR���������������������E�	������Q������-b����\����E���D����R����\�����tƅ�����E��������?���E��M���p���  �EP�MQ�vL�����Ѕ�t�t  ������P��p����p���������������������E�
��|�������|����������ɉ����vej ������P��p�����o���������������������E�   ��|�������|����������m���0�M�wq����;�uǅ���   �
ǅ���    �������Z����E�
   ��|�����t��|������������o���E�   ��|�����t��|�����������o����Z�����t?�M軅��������R��p����o��������������P�M��R���������ho���!  �����Q��p����+c���������������������E���|�������|����������v�����vej ������Q��p�����b���������������������E�   ��|�������|����������3l���0�M�$p����;�uǅ���   �
ǅ���    �������S����E�   ��|�����t��|��������~n���E�   ��|�����t��|����������Zn����S�����tF�M�h�����H���P��p����b��������������Q�M��QQ����H����n��ƅw�����   ��,���R��p����pm���������������;�����uǅ ���   �
ǅ ���    �� �����_�����,����m����_�����t�f������R��p����pa���������������چ����uǅ,���   �
ǅ,���    ��,�����[����������Tm����[�����tƅw�����  ǅT���    ��p���膑����8�����d���R��p����cV���E���d����CS����u3�f��B������p�������f��B���f��B���f��H�����H�����t��d����I��� ��|e��M�˂���MQ�UR��Z��������t?�M��m����Q�UR��x������h�����h���
s��h�������Q�M���H����M  j j�M��>S���E�ǅx���    ��M�L����UR�EP�XZ�����ȅ���   �M�am����R�EP�Xx������h�����h���
sW��h�������R�M��eH����x���P�M���G�����t(��x���R�M��G���������������������
�K��x���P�M��G�����t�M��l������H���;�t�"�j j�M��U����x�������x���������x��� u�.��x���R�M��8G��� ��~��x�������x����ƅ������d����TG����L�������������   ��x��� ��   ��L������u
�   �   ��x�������x���t��L����0��x���Q�M��F���;�u(��x��� u(��L����0��x���Q�M��F���;�}	ƅ�����%�   �� ��L������~��L�������L����A�����������t �E��M��L���E���d����|L����  �E��M��kL����p����1g��f��D����UR�EP�X�����ȅ���   ��D�������   �M�k������D���;���   �UR�M����P��W��������t\��T���;�8���}N�M��j����R�EP��u������h�����h���
s'��h�������R�M���E����T�������T���눋�T���;�8���}ƅ�����M��YO����u	ƅ�����+���T�������T�����T���;�8���}j0�M��sE�����E���d����9K���   ��`���u�vƅo��� ��M��~���MQ�UR��V��������t)�M��i����QjH��$�����V���Ѕ�t	ƅo���븋�`�����4����� u��o�����uƅ������������������  �M�胁������  �������|V���E���,���Q�M���|���������������������E�������P��������O���E���,����lI����M��}����P���Q�M���H����������������|����E���|����� ��|�����|���Q�������Ay�����X���Ѕ�t@�EP�MQ�U�����Ѕ�t)�M�h�����������.y��� ;�uǅ0���   �
ǅ0���    ��0�����]����E�   ��|����� t��|���ߍ�P����H����]�����t������8���Q�M���G���������������������E�������P��������W����g����E���8����8H����g�����tƅ�����E��������5����������tj �M��Sy�����w�����tj-jj �M��܄���M�Q�M�?H����|�����@��|����E��M��H���E������M��f���E�M�d�    Y^�M�3��1Y����]� ��Y���R�����  �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��,8���E��}� t�E�P�M����AB���M�Q��z�����M����n���Ѕ�u�M����G���E���E���E��]�������������������������������U��Q�M��E�� ��]�����������������U����M��E��H�9 t�U��B,��M���E�    �E����]�����������������U����M��E��H�9 t�U��B,��M���E�    �E����]�����������������U����M��E��H,����E��H,��U��B��M��U��B����U��B��E���]��������������������������������U����M��E��H,����E��H,��U��B��M��U��B����U��B��E���]��������������������������������U����M��M��[��;Es�M���p���E��H;Ms�U��BP�MQ�M���7���J�U��t2�}s,�E��M;Hs�U�U��	�E��H�M��U�Rj�M���u����} u
j �M��lZ���} v	�E�   ��E�    �E��]� �����������������������������������������U����M��M���-��;Es�M��b����E��H;Ms�U��BP�MQ�M���R���J�U��t2�}s,�E��M;Hs�U�U��	�E��H�M��U�Rj�M��RQ����} u
j �M��WD���} v	�E�   ��E�    �E��]� �����������������������������������������U����E�ŝ��E� �E�ŝ��E�    �	�E����E��M�;Ms�UU��3E��E�iM�� �M��ԋE���]��������������������������U����E�E��M��%�U����U��E�� t�M��+�U����U��E��t�M��#�U����U��   k� �U�
��Lt�   k� �E��M���E����E��-�M��I�U����U��E�� 6�M����M��U��4�E����E��M��   �M�}�   u�E�o�:�}�   t�   �� �E��M���U��t�E�X��E�x�E��E��M��M��U��E���M����M��U�� �E��]��������������������������������������������������������������������������������������U����E�E��M��%�U����U��E�� t�M��+�U����U��E��t�M��#�U����U��   k� �U�
��Lt�   k� �E��M���E����E��-�M��I�U����U��E�� 6�M����M��U��4�E����E��M��   �M�}�   u�E�o�:�}�   t�   �� �E��M���U��t�E�X��E�x�E��E��M��M��U��E���M����M��U�� �E��]��������������������������������������������������������������������������������������U����M��E��8 t.�M��	�z��f�E��Ma��f�E��U�R�E�P�+�����ȅ�t�U��    �E��@��M��A ��]�������������������������������������U����M��E��8 t.�M��	�k��f�E��v��f�E��U�R�E�P�3q�����ȅ�t�U��    �E��@��M��A ��]�������������������������������������U��j�h��d�    PQ��@���3ŉE�SVWP�E�d�    �e��M��E�P�M��`���}���,�   ���M��b���E��M��A    �U��B    �E��@    �M��A    �E�    �U���,Rj �E��HQ�d:�����E��U��E��B�M�Qj �M��@����M��7Y��j j �c`���K���E�������E������U��B(��t�M��Q(�U��	�E��H)�M��U��E��P�M��y |	�U��z|
�E��@    �M��Q.R�E��H*Q�U��B+P�M��� Q�M��3���U��B/P�M��Q,R�E��H-Q�U���$R�M��}3���E��t,jh ��M��� Q��5����jh ��U���$R�5�����M�d�    Y_^[�M�3��(K����]� �������������������������������������������������������������������������������������������������������������������������U��j�h��d�    PQ��@���3ŉE�SVWP�E�d�    �e��M��E�P�M�^���}���,�   ���M�`���E��M��A    �U��B    �E��@    �M��A    �E�    �U���,Rj �E��HQ�$8�����E��U��E��B�M�Qj �M���C����M��=��j j �#^�������E�������E������U��B(��t�M��Q(�U��	�E��H)�M��U��E��P�M��y |	�U��z|
�E��@    �M��Q.R�E��H*Q�U��B+P�M��� Q�M��r���U��B/P�M��Q,R�E��H-Q�U���$R�M��r���E��t,jh ��M��� Q�3����jh ��U���$R�}3�����M�d�    Y_^[�M�3���H����]� �������������������������������������������������������������������������������������������������������������������������U���4���3ŉE�VW�M̍E�P�M�\���}̃��   ���_^�M�3��-H����]� ������������������������������U���4���3ŉE�VW�M̍E�P�M�3\���}̃��   ���_^�M�3���G����]� ������������������������������U����M��E�P�M�2m����P�E��H�P��]� �����������������������U����M��E�P�M��l����P�E��H�P��]� �����������������������U���D���3ŉE�VW�M̍E�P�M�&���M̃����P�Q�P�Q�@�A�M�Q�M�+[���}̃��   ���_^�M�3���F����]� ��������������������������������������U���D���3ŉE�VW�M̍E�P�M�%���M̃����P�Q�P�Q�@�A�M�Q�M�Z���}̃��   ���_^�M�3��5F����]� ��������������������������������������U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��j�h��d�    PQ��   ���3ŉE�SVWP�E�d�    �e��M��M�p[���E��E�P�M�hY���M��A    �U��B    �E��@    �E�    �M��t	�E��Q�	�U��B�E��M�Q�M�Y����p�����p���Rj �E�P��2������x����M���x����Q�M�o���E��E�Pj �M�Q�$������|����U���|����B�M�',����t����M�Qj ��t���R�S$�����E��E��M��H��M��EF��j j �zX���4 ��E�������E������U��t0�E�Pj j.�N@�����M�f�A�U�Rj j,�7@�����M�f�A���,�   �u����U�Rj �M��W���M�d�    Y_^[�M�3��C����]� ������������������������������������������������������������������������������������������������������������������U��j�h0�d�    PQ��   ���3ŉE�SVWP�E�d�    �e��M��M�@Y���E��E�P�M�8W���M��A    �U��B    �E��@    �E�    �M��t	�E��Q�	�U��B�E��M�Q�M��V����p�����p���Rj �E�P�0������x����M���x����Q�M�Vm���E��E�Pj �M�Q�f������|����U���|����B�M��)����t����M�Qj ��t���R�Rf�����E��E��M��H��M��`��j j �JV���d��E�������E������U��t0�E�Pj j.�q�����M�f�A�U�Rj j,�jq�����M�f�A���,�   �u����U�Rj �M��8%���M�d�    Y_^[�M�3��A����]� ������������������������������������������������������������������������������������������������������������������U��j�hp�d�    PQ��SVW���3�P�E�d�    �e��M�E��@    �M��A    �U��B    �E�    �EPj �M��	M���M�l���E�M�U�Q��M��Ya��j j ��T������E�������E������M�d�    Y_^[��]� ���������������������������������������������U��j�h��d�    PQ��SVW���3�P�E�d�    �e��M�E��@    �M��A    �U��B    �E�    �EPj �M�� ���M�9k���E�M�U�Q��M���/��j j ��S������E�������E������M�d�    Y_^[��]� ���������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M�E�P�M�H���E��M��M��E�    �U�R�M���@,���E������M��Ug���M�d�    Y��]� �����������������������������U��j�h�d�    P�����3�P�E�d�    �M�E�P�M�G���E��M��M��E�    �U�R�M���+���E������M���f���M�d�    Y��]� �����������������������������U��Q�M��} t#�M��W2��9Er�M��J2���M��Q�P;Ew2������]� ������������������U��Q�M��} t#�M���N��9Er�M���N���M��Q�P;Ew2������]� ������������������U��j�hP�d�    P��   ���3ŉE�P�E�d�    h�  h���EP�w*�����}$ v�M ���+t�E ���-u	�E�   ��E�    �U��U��M�Bc��%   =   u@�E���;E$w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M��U�R�M�A����|�����|�����t����E�    ��t���Q�qM�����E��E������M��5��j �U$R�M��,���E�   j �M���0��P�E E$P�   k� U R�M��!\���E�P�M��@����x�����x����M��E��U�R�EG�����E��E��M������E�P�M��c=���E�j �M��+&���E��M����tz�E����~p�M��S��f�E��U����tY�M����~O�E���U$+U�;�s?�E���U$+щU$�E�Pj�M$Q�M��O���   �� �E����~	�U����U�뜍M��;g���E$�M��F���E��U��}� |%�}� v�M��F��;E$v�M�F��+E$�E���E�    �E��E��M�@a��%�  �E��}�@ty�}�   tp�M�Q�UR�EP�MQ��T���R�EP�8h������P�M�U�E�    �E�Pj �M��S/��P�MQ�UR��l���P�MQ��E������@�U�E�   �}�   um�M�Qj �M��/��P�UR�EP��D���Q�UR�E������P�M�U�E�P�MQ�UR�EP��\���Q�UR�g������P�M�U�E�    �5�E�Pj �M��.��P�MQ�UR��L���P�MQ�-E������@�U�E�M$+M�Q�U�R�M��i.��P�EP�MQ��d���R�EP��D������P�M�Uj j �M��*���E�P�MQ�UR�EP�MQ�UR��f�����E��M��(���E������M��)���E�M�d�    Y�M�3��@9����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��   ���3ŉE�P�E�d�    h�  h���EP�a�����}$ v�M ���+t�E ���-u	�E�   ��E�    �U��U��M��]��%   =   u@�E���;E$w5�M M����0u'�E E��H��xt�U U��B��Xu	�M����M��U�R�M�<����|�����|�����t����E�    ��t���Q�t�����E��E������M�����j �U$R�M��xY���E�   j �M��%A��P�E E$P�   k� U R�M��(���E�P�M�;����x�����x����M��E��U�R�������E��E��M��`���E�P�M��)0���E�j �M��� ���E��M����tz�E����~p�M��;��f�E��U����tY�M����~O�E���U$+U�;�s?�E���U$+щU$�E�Pj�M$Q�M��@���   �� �E����~	�U����U�뜍M��\���E$�M�A���E��U��}� |%�}� v�M�fA��;E$v�M�YA��+E$�E���E�    �E��E��M��[��%�  �E��}�@ty�}�   tp�M�Q�UR�EP�MQ��T���R�EP�=S������P�M�U�E�    �E�Pj �M��y?��P�MQ�UR��l���P�MQ�>������@�U�E�   �}�   um�M�Qj �M��6?��P�UR�EP��D���Q�UR�U>������P�M�U�E�P�MQ�UR�EP��\���Q�UR�R������P�M�U�E�    �5�E�Pj �M���>��P�MQ�UR��L���P�MQ��=������@�U�E�M$+M�Q�U�R�M��>��P�EP�MQ��d���R�EP�=������P�M�Uj j �M�%���E�P�MQ�UR�EP�MQ�UR��Q�����E��M��;#���E������M���@���E�M�d�    Y�M�3���3����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hL�d�    P���   ���3�P�E�d�    j j �$�����   ������#Uu�   �} um��G���E�jUh��E�PjD�e#�����E��E�    �}� tj �MQ�M��mT���E���E�    �U�U��E������������P�E�P�M��*��� ������P�MQ��B����P�M�*��j j �aA�����   ������#Uu�   �} uy�GG����P���jVh���P���Pj�"�����E��E�   �}� tj �MQ�M��V���E���E�    �U���x����E�����������P��x���P�M�*��� �������P�MQ��/����P�M��)��j j ������   ������#Uu�   �} uy�F����8���jWh���8���Pj��!�����E��E�   �}� tj �MQ�M��w`���E���E�    �U؉�p����E���������V��P��p���P�M�K)��� ����:��P�MQ�����P�M�))��j j ��(�����   ������#Uu�   �} u{��E����H���jXh���H���Pj�+!�����E��E�   �}� tj j �MQ�M��.���E���E�    �UЉ�h����E�����������P��h���P�M�(��� ����x��P�MQ��:����P�M�g(��j j ��2�����   ������#Uu�   �} uy�E����(���jYh���(���Pj�i �����E��E�   �}� tj �MQ�M��*H���E���E�    �Uȉ�`����E������������P��`���P�M��'��� ������P�MQ�`>����P�M�'��j j �N�����   ������#Uu�   �} uy�ED����@���jZh���@���Pj������E��E�   �}� tj �MQ�M���(���E���E�    �U���X����E�����������P��X���P�M�	'��� �������P�MQ��J����P�M��&��j j �5>�����   ������#Uu�   �} us�C����0���j[h���0���Pj�������E��E�   �}� tj �MQ�M��~E���E���E�    �U�U��E���������W��P�E�P�M�O&��� ����>��P�MQ��!����P�M�-&��j j �G5�����   ������#Uu�   �} uy��B����|���j\h���|���Pj�/�����E��E�   �}� tj �MQ�M��;���E���E�    �U܉�t����E�����������P��t���P�M�%��� ����~��P�MQ�8����P�M�m%��j j �G�����   ������#Uu�   �} u{�B����l���j]h���l���PjX�o�����E��E�   �}� tj j �MQ�M��Y���E���E�    �Ủ�d����E������������P��d���P�M��$��� ������P�MQ�P����P�M�$��j j ��\�����   ������#Uu�   �} u{�IA����\���j^h���\���PjX������E��E�	   �}� tj j �MQ�M��J���E���E�    �U���T����E�����������P��T���P�M�$��� �������P�MQ�p+����P�M��#��j j �*�����   ������#Uu�   �} uy�@����L���j_h���L���PjD�������E��E�
   �}� tj �MQ�M��0���E���E�    �U���D����E���������V��P��D���P�M�K#��� ����:��P�MQ�4����P�M�)#��j j �c�����   ������#Uu�   �} uy��?����<���j`h���<���Pj�+�����E��E�   �}� tj �MQ�M��B���E���E�    �U���4����E�����������P��4���P�M�"��� ����z��P�MQ�D����P�M�i"��j j ��)�����   ������#Uu�   �} uy�?����,���jbh���,���Pj4�k�����E��E�   �}� tj �MQ�M���M���E���E�    �U���$����E������������P��$���P�M��!��� ������P�MQ�Y����P�M�!���M�d�    Y��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h,�d�    P���   ���3�P�E�d�    j j �?#�����   ������#Uu�   �} um�;���E�j-h��E�PjD�������E��E�    �}� tj �MQ�M��(���E���E�    �U�U��E���������c��P�E�P�M�[��� ����J��P�MQ������P�M�9��j j �PD�����   ������#Uu�   �} uy��:����P���j.h���P���Pj�;�����E��E�   �}� tj �MQ�M��S���E���E�    �U���x����E������x����P��x���P�M���� �x����P�MQ�����P�M�y��j j �[�����   ������#Uu�   �} uy�:����8���j/h���8���Pj�{�����E��E�   �}� tj �MQ�M�����E���E�    �U؉�p����E������|�����P��p���P�M����� �|�����P�MQ��B����P�M���j j �&$�����   ������#Uu�   �} u{�W9����H���j0h���H���Pj������E��E�   �}� tj j �MQ�M��G���E���E�    �UЉ�h����E������t��$��P��h���P�M���� �t����P�MQ�����P�M����j j ������   ������#Uu�   �} uy�8����(���j1h���(���Pj�������E��E�   �}� tj �MQ�M��N���E���E�    �Uȉ�`����E���������d��P��`���P�M�Y��� ����H��P�MQ�N����P�M�7��j j �$�����   ������#Uu�   �} uy��7����@���j2h���@���Pj�9�����E��E�   �}� tj �MQ�M��1���E���E�    �U���X����E�����������P��X���P�M���� ������P�MQ�Q$����P�M�w��j j ��������   ������#Uu�   �} us�7����0���j3h���0���Pj�y�����E��E�   �}� tj �MQ�M��Z3���E���E�    �U�U��E����������
��P�E�P�M����� �����
��P�MQ������P�M���j j ��������   ������#Uu�   �} uy�[6����|���j4h���|���Pj������E��E�   �}� tj �MQ�M������E���E�    �U܉�t����E���������*
��P��t���P�M���� ����
��P�MQ�p�����P�M����j j �#�����   ������#Uu�   �} u{�5����l���j5h���l���PjX�������E��E�   �}� tj j �MQ�M��A���E���E�    �Ủ�d����E���������h	��P��d���P�M�]��� ����L	��P�MQ�����P�M�;��j j �������   ������#Uu�   �} u{��4����\���j6h���\���PjX�=�����E��E�	   �}� tj j �MQ�M��QB���E���E�    �U���T����E�����������P��T���P�M���� ������P�MQ�UB����P�M�y��j j �#�����   ������#Uu�   �} uy�4����L���j7h���L���PjD�{�����E��E�
   �}� tj �MQ�M�����E���E�    �U���D����E������������P��D���P�M����� �������P�MQ�.N����P�M���j j ��8�����   ������#Uu�   �} uy�W3����<���j8h���<���Pj������E��E�   �}� tj �MQ�M������E���E�    �U���4����E������t��&��P��4���P�M���� �t��
��P�MQ�����P�M����j j �^ �����   ������#Uu�   �} uy�2����,���j:h���,���Pj4�������E��E�   �}� tj �MQ�M��^H���E���E�    �U���$����E���������f��P��$���P�M�[��� ����J��P�MQ�����P�M�9���M�d�    Y��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EP��$�������E�jAh���K/��P3ɋE��   �������Q��������E�E�E��M�Q�UR�E�P�8�����E���]����������������������������U����M��E��H(��u,�}w&�}w �}wkU�E��kU(�����E���E� ��M��M�j�U�Rj�EP�<������]� �������������������������U����M��E��H(��u,�}w&�}w �}wkU�E��kU(�����E���E� ��M��M�j�U�Rj�EP�������]� �������������������������U����M��E��xr�M��QR������E��	�E����E��E���]���������������������������U����M��E��xr�M��QR�M�����E��	�E����E��E���]���������������������������U����M��E��xr�M��QR������E��	�E����E��E���]���������������������������U����M��E��xr�M��QR�������E��	�E����E��E���]���������������������������U��j�h��d�    P�����3�P�E�d�    �E�   �} u	�E�    ��EP�M��;���E��M��M��E� �M�����E������M�����E�M�d�    Y��]������������������������������������U��j�h �d�    P�����3�P�E�d�    �E�   �} u	�E�    ��EP�M��5���E��M��M��E� �M������E������M������E�M�d�    Y��]������������������������������������U����M�E�8 t.�M�	���f�E��M)��f�E��U�R�E�P�������ȅ�t�U��    ��E�P��0�����M�f�A�U��B�E�f�@��]����������������������������������U����M�E�8 t.�M�	�E	��f�E��>��f�E��U�R�E�P�#9�����ȅ�t�U��    ��E�P�D"�����M�f�A�U��B�E�f�@��]����������������������������������U����M��E��H �9 t�U��B0��M���E�    �E����]�����������������U����M��E��H �9 t�U��B0��M���E�    �E����]�����������������U����M��E��H0����E��H0��U��B ��M��U��B ����U��B ��E���]��������������������������������U����M��E��H0����E��H0��U��B ��M��U��B ����U��B ��E���]��������������������������������U��j�h8�d�    P���3�P�E�d�    �E�    ��E ���E �M�;���M�*���}  v �M�X��f���R�M������#�����E�M��U�P�E������M�S����E�M�d�    Y��]����������������������������������������U��j�hh�d�    P���3�P�E�d�    �E�    ��E ���E �M�����M�1���}  v �M�+1��f���R�M������_�����E�M��U�P�E������M�����E�M�d�    Y��]����������������������������������������U����E���E�M�>:���M���M�} v�U�P�M������E"���ȋM�U��E�A�E]���������������������������������U����E���E�M������M���M�} v�U�P�M�
�����\���ȋM�U��E�A�E]���������������������������������U��j�h)�d�    P��  ���3ŉE�P�E�d�    ��X����E�    h  h(��EP�
������M��tK������R�M����������������������E�������Q��������8����E� �������C����I��t���R�M�B����������������|����E���|���Q��4������8����E� ��t���������U�R��8����!���E���8���������������� }������؉����������������������@����M$��;��;�@���w(�E@P�M$�;����@���+ȃ�Qj �M$��#����   �M�����������   �M������ ����   ��8������f������M�������0����M$�A;��+�@�����(�����0������tx��0������~k��0����;�(���sZ��0������(���+�(��������Qj��(���R�M$�#���   �� ��0������~��0�������0����z����M��=���E��M ��tH��`���R��8��������� �� ����M�Q��8����X����x�����x���R�M��� ���M�������L��H���P��8����
������ �����H���R��8�������������������P�M�� ����H����u����M���<���E��M�I4����t2��d���Q��8����*��������������R�M��V ����d����*���ƅ?��� ǅD���    ǅ4���    ���4�������4�����4����  ��4����� �����,�����,����� ��,�����,���X��   ��,�����0?�$�?�M��79���D�����D����   �M��9���D�����D����   ��@��� vǅ���   �
ǅ���    �M$��8��;�@���w�M$��8����@���+ȃ�������
ǅ���    �M$�8�����������D�����D������D�������D�����4���tƅ?���������M��������������������� |1	������ v&�M����;�D���v�M����+�D���������
ǅ���    �������D����M�]2��%�  ����������@tO�����   u��?�����u8��D���R�EP�MQ�UR������P�������P�M�UǅD���    ǅ4���    ���4�������4�����4����  ��4����� �����$�����$����� ��$�����$���X��  ��$������?�$��?�M��07��P�����P�M��7����������������������E����̉�@���������R�9����8����EP�MQ������R�;������������������P�M�U�E������������5  �M��6������   j��$���P�M������������������������E����̉�0���������R�y8����L����EP�MQ������R�l:������������������P�M�U�E���$����B����  ��@��� ��   �M$� 6��P�����P�M$�����������������������E����̉�P���������R��7����p����EP�MQ������R��9������������������P�M�U�E�����������  �M$�s5��;�@����	  �E@Pj �M��������V����������8����{:����Qj �M�������/��������M$�5����@���+�R�E@P�MQ�UR��|���P�M�������P�M�U�M$��4��P������P�M$������������������������E�	���̉�d���������R��6����<����EP�MQ��l���R�8������������������P�M�U�E������������y  �M$�V4��+�@���P������P�M$�W����������������������E�
���̉�\���������R�/6����D����EP�MQ��t���R�"8������������������P�M�U�E��������������8����9����Pj �M� �����������B����@���Q��@���R������P������Q�M$�����������������������E��������3���������������������E����̉�T���������R�S5����4����EP�MQ������R�F7������������������P�M�U�E������������E������������mj�EP�MQ�UR������P��������P�M�U�����   u8��D���P�MQ�UR�EP������Q���������@�U�EǅD���    ������M��i2������   �M��X2����Pj�� ���Q������R�M��S����������������� ����E��� ����A���������������������E����̉�l���������R�
4����h����EP�MQ������R��5������������������P�M�U�E��� ���������E������������j j �M������D���P�MQ�UR�EP�MQ��������E��M�������E��M�������E� �M������E������M$�����E�M�d�    Y�M�3��G����]�< �7�67*7�7�7 �I T=�8�9":}=�= ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h)�d�    P��  ���3ŉE�P�E�d�    ��X����E�    h  h(��EP�x*�����M��tK������R�M����������������������E�������Q�.$������8����E� �������C����I��t���R�M�B����������������|����E���|���Q�K�������8����E� ��t���������U�R��8����N����E���8����J1������������ }������؉����������������������@����M$�&��;�@���w(�E@P�M$��%����@���+ȃ�Qj �M$�������   �M�����������   �M������ ����   ��8����o$��f������M�������0����M$�%��+�@�����(�����0������tx��0������~k��0����;�(���sZ��0������(���+�(��������Qj��(���R�M$�����   �� ��0������~��0�������0����z����M������E��M ��tH��`���R��8�������� �� ����M�Q��8����9�����x�����x���R�M��{����M��B���L��H���P��8����������� �����H���R��8����
��������������P�M��0�����H�����
���M��:���E��M�I$����t2��d���Q��8��������������������R�M��������d����
��ƅ?��� ǅD���    ǅ4���    ���4�������4�����4����  ��4����� �����,�����,����� ��,�����,���X��   ��,�����0O�$�O�M��y#���D�����D����   �M��`#���D�����D����   ��@��� vǅ���   �
ǅ���    �M$�(#��;�@���w�M$�#����@���+ȃ�������
ǅ���    �M$��"�����������D�����D������D�������D�����4���tƅ?���������M��������������������� |1	������ v&�M����;�D���v�M����+�D���������
ǅ���    �������D����M�]"��%�  ����������@tO�����   u��?�����u8��D���R�EP�MQ�UR������P�r�������P�M�UǅD���    ǅ4���    ���4�������4�����4����  ��4����� �����$�����$����� ��$�����$���X��  ��$������O�$��O�M��r!��P�����P�M������������������������E����̉�@���������R�)�����8����EP�MQ������R�4������������������P�M�U�E�������9����5  �M��� ������   j��$���P�M��0���������������������E����̉�0���������R������L����EP�MQ������R�������������������P�M�U�E���$��������  ��@��� ��   �M$�B ��P�����P�M$����������������������E����̉�P���������R�������p����EP�MQ������R�������������������P�M�U�E�������	����  �M$���;�@����	  �E@Pj �M��������������j����8����f����Qj �M�������g������C���M$�]����@���+�R�E@P�MQ�UR��|���P��������P�M�U�M$�%��P������P�M$�y���������������������E�	���̉�d���������R�������<����EP�MQ��l���R��������������������P�M�U�E�������������y  �M$���+�@���P������P�M$�����������������������E�
���̉�\���������R�I�����D����EP�MQ��t���R�T������������������P�M�U�E��������Y�����8���������Pj �M�-������������������@���Q��@���R������P������Q�M$�}����������������������E�������������������������������E����̉�T���������R�m�����4����EP�MQ������R�x������������������P�M�U�E��������}����E��������n����mj�EP�MQ�UR������P�~�������P�M�U�����   u8��D���P�MQ�UR�EP������Q�D�������@�U�EǅD���    ������M��������   �M������Pj�� ���Q������R�M������������������� ����E��� ��������������������������E����̉�l���������R�$�����h����EP�MQ������R�/������������������P�M�U�E��� ����4����E��������%���j j �M������D���P�MQ�UR�EP�MQ�)������E��M��Q���E��M��E���E� �M������E������M$�*���E�M�d�    Y�M�3��G�����]�< �G�FG*G�G�G �I TM�H�I"J}M�M ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E���E�M�^���} v�MQ�M��������p���ӋU�E��M�J�E]����������������������������U����E���E�M�,����} v�MQ�M�����������ӋU�E��M�J�E]����������������������������U����E���E�M����} v�MQ�M�#������ ���ӋU�E��M�J�E]����������������������������U����E���E�M�l����} v�MQ�M�������������ӋU�E��M�J�E]����������������������������U��Q�M��E��HQ�g������U��BP�X������M��QR�I������E��HQ�:�������]��������������������������U��Q�M��E��HQ�������U��BP��������M��QR��������E��HQ���������]��������������������������U����M��E��u�s�M��yrj�U��B�E�M���Q�U�R�M��C���������} v �EP�M�Q�������P�U���R�������E��H��Q�U�R�E�P�M�������������M��A   �UR�M��h�����]� ����������������������������������������������U����M��E��u�s�M��yrj�U��B�E�M���Q�U�R�M��u������t���} v �EP�M�Q�2�����P�U���R�'������E��H��Q�U�R�E�P�M��.����������M��A   �UR�M��S�����]� ����������������������������������������������U��Q�M��E��HQ�������U��BP��������M��QR���������]�������������������������U��Q�M��E��HQ�������U��BP�������M��QR��������]�������������������������U��Q�M��E��HQ�g������U��BP�X������M��QR�I�������]�������������������������U��Q�M��E��HQ�������U��BP�������M��QR���������]�������������������������U����M�����E��}� t�E�P�M��������M�Q�1�����M���� ���Ѕ�u�M����&����E���E����E��]�������������������������������U����M�� ����E��}� t�E�P�M����-����M�Q������M����
���Ѕ�u�M��������E���E��E��]�������������������������������U����M��E�    �}���P�M�H����E����E��E��]� ����������������U��Q�M�h\[������]������������U��Q�M�h\[�����]������������U��Q�M�hp[�>�����]������������U��Q�M�hp[������]������������U��Q�M��EP�M�������]� �������U��Q�M��EP�M��c�����]� �������U��Q�M�j �EP�u������]� ���������������������U��Q�M�j �EP�N�������]� ���������������������U��Q�M����Pj �MQ�M��"
����]� ���������������U����M��M�F��;Es�M������M�1��+E�E��E�;Es�M��M�U����+B;Ew�M��O���} vZ�M��QU�U�j �E�P�M��2���ȅ�t9�UR�M�
����M�HR�M��(����M��Q�PP�Q������M�Q�M�������E���]� �����������������������������������������������������U����M��E����+H;Mw�M�����} vE�U��BE�E�j �M�Q�M��r���Ѕ�t$�EP�MQ�U��BP�M�������M�Q�M��7����E���]� ������������������������������������������U��Q�M��ĊPj �MQ�M��=�����]� ���������������U����M��M����;Es�M������M���+E�E��E�;Es�M��M�U��Ċ+B;Ew�M������} vZ�M��QU�U�j �E�P�M��+����ȅ�t9�UR�M������M�HR�M��7����M��Q�PP�������M�Q�M�������E���]� �����������������������������������������������������U����M��E��Ċ+H;Mw�M�����} vE�U��BE�E�j �M�Q�M��k����Ѕ�t$�EP�MQ�U��BP�M�������M�Q�M��2����E���]� ������������������������������������������U����M��E�;Eu�a�M�Q�M�����P�U�R�M������P�k���������t�M�yr�UR�M�������!j j�M��3	���EP�:����P�M������E���]� �����������������������������������U��Q�M����Pj �MQ�M�� ����]� ���������������U����M��M�&��;Es�M������M���+E�E��E;E�s�M�M��U�;Uu�EE�P�M������MQj �M�������Ej �U�R�M��������t0�M�Q�M������U�PP�M�����P�=������M�Q�M�������E���]� �������������������������������������������������U��Q�M��E;��u�M����j �MQ�M��|���Ѕ�t�EP�MQj �M�������UR�M��F����E���]� �������������������������U��Q�M�h�  hXo�EP��������MQ�������P�UR�M�������]� ��������������������U��Q�M��} th  hXo�EP�������MQ�M���
���Ѕ�t"�EP�M������M+���Q�U�R�M�����=j �EP�M��~���ȅ�t%�UR�EP�M�����P�������MQ�M��B����E���]� �����������������������������������������������������U����M��E�;Eu�a�M�Q�M����P�U�R�M�����P�J��������t�M�yr�UR�M��X����!j j�M��I����EP������P�M�������E���]� �����������������������������������U��Q�M��ĊPj �MQ�M��������]� ���������������U����M��M�(��;Es�M�������M���+E�E��E;E�s�M�M��U�;Uu�EE�P�M��+���MQj �M������Ej �U�R�M���������t0�M�Q�M�@����U�PP�M�����P��������M�Q�M��I����E���]� �������������������������������������������������U��Q�M��E;Ċu�M����j �MQ�M�������Ѕ�t�EP�MQj �M������UR�M�������E���]� �������������������������U��Q�M�h�  hXo�EP�������MQ������P�UR�M��E�����]� ��������������������U��Q�M��} th  hXo�EP�������MQ�M������Ѕ�t"�EP�M��I����M+���Q�U�R�M�������=j �EP�M�������ȅ�t%�UR�EP�M�����P�f������MQ�M������E���]� �����������������������������������������������������U��EP�MQ�UR�S�����]�������U��E�Mf�f�]����������������U��EP�MQ�UR������]�������U��E�Mf�f�]����������������U��Q�M��E�P�M��Y���P�M����E��]� �����������U��Q�M��E�P�M������P�M�v����E��]� �����������U��Q�M��M��������]��������������U��Q�M��M��C�����]��������������U��Q�} u�E�E���MQ�UR�EP�o������E��E���]�����������������U��Q�} u�E�E���MQ�UR�EP�/������E��E���]�����������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M��EP�MQ�M��R����]� �������������������U��Q�M��EP�MQ�M��=�����]� �������������������U��Q�M��EP�m������]� �������U��Q�M��EP�M������]� �������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M�2���]����U��Q�M�2���]����U��Q�M���]� ���U��Q�M���]� ���U����M�j_h���EP�MQ�>�����j`h���UR�EP�'������M���Q�UR�EP�MQ�UR�c������E��}� }	�E�������}� u	�E�    ��E�   �E��E�E��]� �����������������������������������U����M�j_h���EP�MQ�7�����j`h���UR�EP� ������M���Q�UR�EP�MQ�UR�������E��}� }	�E�������}� u	�E�    ��E�   �E��E�E��]� �����������������������������������U����M��E�    �E��HQ�M�����U����U��E��]� ���������������U����M��E�    �E��HQ�M�����U����U��E��]� ���������������U��Q�M��E��@��]����������������U��Q�M��E��@��]����������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M�3���]����U��Q�M�3���]����U����M��E�    �E��HQ�M�!����U����U��E��]� ���������������U����M��E�    �E��HQ�M�����U����U��E��]� ���������������U��Q�M��E��@��]����������������U��Q�M��E��@��]����������������U����M��E�    �EP�M������M����M��E��]� ������������������U����M��E�    �EP�M������M����M��E��]� ������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M��d���E�    �EP�MQ��������Ѕ�t�E$����U$�
�M��w�����u�E$����U$�
�P�M��p����E��E�    �E�Pj �M�Q�U�R�������]��E�;E�t�}� t�M$����E$���M(�E���U�E��M�J�E������M������E�M�d�    Y�M�3��������]�$ �����������������������������������������������������������������������������������U��j�h��d�    P��H���3ŉE�VP�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M�������E�    �M��*����E��EP�MQ�������Ѕ�t�E$����U$�
�}� u�E$����U$�
�   �E�    �E�P�M(�t���j �M�蜾�����-u+�U��U��E�P�M(�I����   k�
f�L�f��U����U��	�E����E��M�;M�s(�U�R�M��J����0�E�P�M(����f��ux���f��ǋU�E��M�J�E������M��j����E�M�d�    Y^�M�3�������]�$ ����������������������������������������������������������������������������������������������U��j�h�d�    P��P���3ŉE�P�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M��A ���E�    �EP�MQ�ռ�����Ѕ�t�E$����U$�
�M��G�����u�E$����U$�
�P�M��@����E��E�    �E�Pj �M�Q�U�R�O������]��E�;E�t�}� t�M$����E$���M(�E���U�E��M�J�E������M�������E�M�d�    Y�M�3�������]�$ �����������������������������������������������������������������������������������U��j�hX�d�    P��H���3ŉE�VP�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M�������E�    �M�������E��EP�MQ�Y������Ѕ�t�E$����U$�
�}� u�E$����U$�
�   �E�    �E�P�M(����j �M��l������-u+�U��U��E�P�M(�����   k�
f�L�f��U����U��	�E����E��M�;M�s(�U�R�M������0�E�P�M(�X���f��ux���f��ǋU�E��M�J�E������M��:����E�M�d�    Y^�M�3��������]�$ ����������������������������������������������������������������������������������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP�.������E�    �M�Q�M������E��U��U��E�    �E�P�M�A���P�MQ�UR�E�P�M�Q��������E��E������M�蛮���   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R�������E̍EP�MQ�������Ѕ�t�E ����U �
�E�;E�t�}� u	�}���  v�M ����E ��,�   k� �DЃ�-u
3�+M̉M���ỦUċE$f�M�f��U�E��M�J�E�M�d�    Y�M�3�������]�  ������������������������������������������������������������������������������������������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP�>������E�    �M�Q�M�����E��U��U��E�    �E�P�M�Q���P�MQ�UR�E�P�M�Q��������E��E������M�諬���   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R�!������E̍EP�MQ�������Ѕ�t�E ����U �
�E�;E�t�}� u�}��v�M ����E ��*�   k� �DЃ�-u
3�+M̉M���ỦUċE$�Mĉ�U�E��M�J�E�M�d�    Y�M�3�������]�  �����������������������������������������������������������������������������������������������������������U��j�h�d�    P��@���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP�N������E�    �M�Q�U�R�M�����E��E��E��E�    �M�Q�M�]���P�UR�EP�M�Q�U�R�������P�E�P�M�Q�������E��E������M�親���UR�EP�S������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3��~�����]�  �������������������������������������������������������������������������������U��j�hX�d�    P��@���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP��������E�    �M�Q�U�R�M�����E��E��E��E�    �M�Q�M�����P�UR�EP�M�Q�U�R�f�����P�E�P�M�Q��������E��E������M��&����UR�EP��������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3��������]�  �������������������������������������������������������������������������������U���T���3ŉE��M�h)  h���EP�MQ�UR�EP�f������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q������P�U�R�E�P�E������]��}� t�M���QQ�E��$�<������]��UR�EP�u������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3�������]�  ����������������������������������������������������������������������������U���X���3ŉE��M�hA  h���EP�MQ�UR�EP�������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q�?�����P�U�R�E�P��������]��}� t�M���Q���E��$�F������]��UR�EP�#������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��Y�����]�  ��������������������������������������������������������������������������U���X���3ŉE��M�hY  h���EP�MQ�UR�EP��������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q�������P�U�R�E�P��������]��}� t�M���Q���E��$��������]��UR�EP��������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��	�����]�  ��������������������������������������������������������������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�hq  h���EP�MQ�UR�EP�^������E�    �M�Q�M�"����E��U��U��E�    �E�Ph   �MQ�UR�E�P�M�Q��������E��E������M��ϣ���   ��t"�E�P�M�Q�U�R�E�P�b�����3ɉE��M���U�R�E�P�M�Q�U�R� ������E��U��E��E��M��M��UR�EP�'������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E��M$��U�E��M�J�E�M�d�    Y�M�3��R�����]�  ���������������������������������������������������������������������������������������������������U��j�h��d�    P��D���3ŉE�P�E�d�    �M�h   h���EP�MQ�UR�EP�������E�    �M�Q�U�R�M�N����E��E��E��E�    �M�Q�M����P�UR�EP�M�Q�U�R�&�����P�E�P�M�Q�������E��U��E������M������UR�EP�������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3�������]�  ��������������������������������������������������������������������������������������U��j�h�d�    P��D���3ŉE�P�E�d�    �M�h  h���EP�MQ�UR�EP��������E�    �M�Q�U�R�M�����E��E��E��E�    �M�Q�M����P�UR�EP�M�Q�U�R薽����P�E�P�M�Q��������E��U��E������M��S����UR�EP� ������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3��%�����]�  ��������������������������������������������������������������������������������������U��j�h��d�    P��   ���3ŉE�P�E�d�    ��L���h�  h���EP�MQ�UR�EP�h�����ǅx��������M����% @  �'  ��H���Q�M������\�����\�����P����E�    ��P���P�Q�������p����E�������H����Þ��j j�M�輞���E�   ��|���Q��p����G�����@�����@�����8����E���8���P�M������E���|��������j �M������M�Q��p����!�����d�����d�����<����E���<���P�M��W����E��M�賰���M��Z���Pj�MQ�UR��������x����E������M�胰���   ǅh���    ��h���P��`���Q�M�������T�����T�����D����E�   ��D���P�M����P�MQ�UR�E�P��L���Q褺����P��X���R�E�P�'�������l����E�������`����[����M�9�X���t��h��� u��l���w��l�����x����EP�MQ��������Ѕ�t�E ����U �
��x��� }�E ����U �
�*��x��� tǅt���   �
ǅt���    �E$��t�����U�E��M�J�E�M�d�    Y�M�3�������]�  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP�x������E�    �M�Q�M�����E��U��U��E�    �E�P�M�����P�MQ�UR�E�P�M�Q��������E��E������M��;����   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R�������E̍EP�MQ谥�����Ѕ�t�E ����U �
�E�;E�t�}� u	�}���  v�M ����E ��,�   k� �DЃ�-u
3�+M̉M���ỦUċE$f�M�f��U�E��M�J�E�M�d�    Y�M�3�襼����]�  ������������������������������������������������������������������������������������������������������U��j�h�d�    P��P���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP�������E�    �M�Q�M�����E��U��U��E�    �E�P�M�����P�MQ�UR�E�P�M�Q��������E��E������M��K����   k� �LЃ�-u�UщU���EЉE��M��MȍU�R�E�P�M�Q�U�R��������E̍EP�MQ��������Ѕ�t�E ����U �
�E�;E�t�}� u�}��v�M ����E ��*�   k� �DЃ�-u
3�+M̉M���ỦUċE$�Mĉ�U�E��M�J�E�M�d�    Y�M�3�躺����]�  �����������������������������������������������������������������������������������������������������������U��j�hH�d�    P��@���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP�������E�    �M�Q�U�R�M设���E��E��E��E�    �M�Q�M�����P�UR�EP�M�Q�U�R�
�����P�E�P�M�Q�N������E��E������M��F����UR�EP��������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3�������]�  �������������������������������������������������������������������������������U��j�h��d�    P��@���3ŉE�P�E�d�    �M�h�  h���EP�MQ�UR�EP�������E�    �M�Q�U�R�M�.����E��E��E��E�    �M�Q�M�}���P�UR�EP�M�Q�U�R芻����P�E�P�M�Q�������E��E������M��ƕ���UR�EP�|������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U�E��M�J�E�M�d�    Y�M�3�螷����]�  �������������������������������������������������������������������������������U���T���3ŉE��M�h)  h���EP�MQ�UR�EP�������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q覾����P�U�R�E�P�������]��}� t�M���QQ�E��$�ܼ�����]��UR�EP�������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��K�����]�  ����������������������������������������������������������������������������U���X���3ŉE��M�hA  h���EP�MQ�UR�EP�`������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q�V�����P�U�R�E�P�|������]��}� t�M���Q���E��$�������]��UR�EP�̝�����ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3��������]�  ��������������������������������������������������������������������������U���X���3ŉE��M�hY  h���EP�MQ�UR�EP�������E�    �E�    �M�Q�U�R�EP�MQ�UR�E�P�M�Q������P�U�R�E�P�������]��}� t�M���Q���E��$�v������]��UR�EP�|������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�E���M�U��E�A�E�M�3�詳����]�  ��������������������������������������������������������������������������U��j�h��d�    P��P���3ŉE�P�E�d�    �M�hq  h���EP�MQ�UR�EP�������E�    �M�Q�M�·���E��U��U��E�    �E�Ph   �MQ�UR�E�P�M�Q�"������E��E������M��o����   ��t"�E�P�M�Q�U�R�E�P������3ɉE��M���U�R�E�P�M�Q�U�R�������E��U��E��E��M��M��UR�EP�К�����ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E��M$��U�E��M�J�E�M�d�    Y�M�3�������]�  ���������������������������������������������������������������������������������������������������U��j�h�d�    P��D���3ŉE�P�E�d�    �M�h   h���EP�MQ�UR�EP��������E�    �M�Q�U�R�M�����E��E��E��E�    �M�Q�M�=���P�UR�EP�M�Q�U�R�J�����P�E�P�M�Q�V������E��U��E������M�胎���UR�EP�9������ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3��U�����]�  ��������������������������������������������������������������������������������������U��j�hH�d�    P��D���3ŉE�P�E�d�    �M�h  h���EP�MQ�UR�EP�H������E�    �M�Q�U�R�M�^����E��E��E��E�    �M�Q�M����P�UR�EP�M�Q�U�R躲����P�E�P�M�Q�|������E��U��E������M������UR�EP詗�����ȅ�t�U ����M ��U�9U�t�}� t�E ����U �
��E$�M���U��P�E�M��U�P�E�M�d�    Y�M�3��Ů����]�  ��������������������������������������������������������������������������������������U��j�h��d�    P��   ���3ŉE�P�E�d�    ��L���h�  h���EP�MQ�UR�EP������ǅx��������M�8���% @  �'  ��H���Q�M賲����\�����\�����P����E�    ��P���P��������p����E�������H����c���j j�M������E�   ��|���Q��p���贗����@�����@�����8����E���8���P�M�趢���E���|�������j �M��ƺ���M�Q��p����������d�����d�����<����E���<���P�M��i����E��M��ҹ���M��]���Pj�MQ�UR��������x����E������M�袹���   ǅh���    ��h���P��`���Q�M�{�����T�����T�����D����E�   ��D���P�M����P�MQ�UR�E�P��L���Q�ȯ����P��X���R�E�P�Ǻ������l����E�������`���������M�9�X���t��h��� u��l���w��l�����x����EP�MQ舔�����Ѕ�t�E ����U �
��x��� }�E ����U �
�*��x��� tǅt���   �
ǅt���    �E$��t�����U�E��M�J�E�M�d�    Y�M�3�荫����]�  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��p���3�P�E�d�    �M��E�P�M�^����E܋M܉M��E�    �U�R�\������E��E������M�� ����E�    �E(�E�M��A�M�}�8�K  �U�����$����M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��������P�M�U�  �E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��+�����@�U�E��  h`��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��������P�M�U�  �E�P�M�Qjcj �UR�EP�M�Q�G������U �M ��U ���ukM�d��l  �U$�J�Q  �E�P�M$��Qjj�UR�EP�M�Q��������U �M ��  h|��U$R�E P�MQ�UR�EP�MQ�UR�E�P�M�������P�M�U��  �E�P�M$��Qjj �UR�EP�M�Q茐�����U �M ��  �U�R�E$��Pjj �MQ�UR�E�P�Z������M �U ��~  �E�P�M$��Qhn  j�UR�EP�M�Q�%������U �M ��I  �U�R�E�Pjj�MQ�UR�E�P��������M �U ��E ���u�U���E$�P�  �M�Q�U$��Rj;j �EP�MQ�U�R讏�����M �U ���  h���E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��������@�U�E�  h��j �MQ�UR�P������E�}� }�E ����U �
�kE��M$A�U$�B�Q  h���E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��K�����@�U�E�  h���M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�������P�M�U��  �E�P�M$Qj;j �UR�EP�M�Q脎�����U �M ��  h���U$R�E P�MQ�UR�EP�MQ�UR�E�P�M�������P�M�U�k  �E�P�M$��Qj5j �UR�EP�M�Q�������U �M ��9  �U�R�E$��Pjj �MQ�UR�E�P�������M �U ��  �E�P�M$��Qj5j �UR�EP�M�Q豍�����U �M ���   hБ�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��������P�M�U�   �E�P�M�Qjcj �UR�EP�M�Q�E������U �M ��U ���u �}�E}�M��d�M���U�U��E$�M��H�B�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M�������P�M�U��E ����U �
�EP�MQ�T������Ѕ�t�E ����U �
�E�M��U�P�E�M�d�    Y��]�( �I $�\�њL�����g�W���Ý �d�)�����"���֜�2���Ӟ^� 	
	 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h(�d�    P��p���3�P�E�d�    �M��E�P�M�����E܋M܉M��E�    �U�R�O������E��E������M�����E�    �E(�E�M��A�M�}�8�K  �U������$�$��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�踁����P�M�U�  �E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��,�����@�U�E��  h`��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��������P�M�U�  �E�P�M�Qjcj �UR�EP�M�Q�������U �M ��U ���ukM�d��l  �U$�J�Q  �E�P�M$��Qjj�UR�EP�M�Q�ү�����U �M ��  h|��U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��3�����P�M�U��  �E�P�M$��Qjj �UR�EP�M�Q�c������U �M ��  �U�R�E$��Pjj �MQ�UR�E�P�1������M �U ��~  �E�P�M$��Qhn  j�UR�EP�M�Q��������U �M ��I  �U�R�E�Pjj�MQ�UR�E�P�ͮ�����M �U ��E ���u�U���E$�P�  �M�Q�U$��Rj;j �EP�MQ�U�R腮�����M �U ���  h���E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��������@�U�E�  h��j �MQ�UR�)������E�}� }�E ����U �
�kE��M$A�U$�B�Q  h���E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��e�����@�U�E�  h���M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��(�����P�M�U��  �E�P�M$Qj;j �UR�EP�M�Q�[������U �M ��  h���U$R�E P�MQ�UR�EP�MQ�UR�E�P�M�������P�M�U�k  �E�P�M$��Qj5j �UR�EP�M�Q�������U �M ��9  �U�R�E$��Pjj �MQ�UR�E�P躬�����M �U ��  �E�P�M$��Qj5j �UR�EP�M�Q般�����U �M ���   hБ�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��������P�M�U�   �E�P�M�Qjcj �UR�EP�M�Q�������U �M ��U ���u �}�E}�M��d�M���U�U��E$�M��H�B�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M�������P�M�U��E ����U �
�EP�MQ�������Ѕ�t�E ����U �
�E�M��U�P�E�M�d�    Y��]�( �I ��̢A�����+�פǥ�3�p�Ԧ�����]���	�F������C�Χ 	
	 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hX�d�    P��D���3�P�E�d�    �M�h  h��EP�MQ�UR�EP������h  h��M$Q�������U�R�M�F����E��E��E��E�    �M�Q�D������E��E������M��w���M��'����E�}� u�E�   �UR�EP蝞�����ȅ�t�  �M�(�����Rj�M�蓿������u?�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��,�����P�M�U�E�   �   �}�u>�E�P�M$��Qjj�UR�EP�M�Q�u������U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P�1������M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M���~����@�U�E�MQ�UR�@���������t'�M�	�����QjH�M��t����Ѕ�t
�M脤���EP�MQ�������Ѕ�t<j �M�ɑ����P�M��e����E��M��:t�U��,t	�E��/u�M�/����MQ�UR����������t'�M�x�����QjH�M������Ѕ�t
�M�����EP�MQ誜�����Ѕ�t��   �M�5�����Pj�M�蠽���ȅ�uW�}�u�U ����M ��@�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��$�����P�M�U�}�u�E�   �w�}�t�}�u>�E�P�M$��Qjj�UR�EP�M�Q�d~�����U �M ��U$�B���M$�A�-�U�R�E$��Pjj�MQ�UR�E�P�&~�����M �U ��EP�MQ�j������Ѕ�t'�M�3�����PjH�M�螼���ȅ�t
�M订���UR�EP�,������ȅ�t<j �M������R�M�菒���E��E��:t�M��,t	�U��/u�M�Y����EP�MQ�ٿ�����Ѕ�t'�M袏����PjH�M������ȅ�t
�M�����UR�EP�Ԛ�����ȅ�t�U ����M ��  �M�R�����Rj�M�轻������uM�}�t�M ����E ��3�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��A�����P�M�U�   �}�u>�E�P�M$��Qjj�UR�EP�M�Q�|�����U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P�M|�����M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��{����@�U�E�MQ�UR蕙��������t�M ����E ��M�U��E�A�E�M�d�    Y��]�  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��D���3�P�E�d�    �M�h  h��EP�MQ�UR�EP軨����h  h��M$Q�:������U�R�M�Ɩ���E��E��E��E�    �M�Q�'r�����E��E������M��o���M��q���E�}� u�E�   �UR�EP�&z�����ȅ�t�  �M跟����Rj�M��Ќ������u?�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�������P�M�U�E�   �   �}�u>�E�P�M$��Qjj�UR�EP�M�Q�<������U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P��������M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�������@�U�E�MQ�UR苋��������t'�M蘞����QjH�M�豋���Ѕ�t
�M�C����EP�MQ�M������Ѕ�t<j �M�X�����P�M��;s���E��M��:t�U��,t	�E��/u�M�����MQ�UR�����������t'�M������QjH�M�� ����Ѕ�t
�M貲���EP�MQ�3x�����Ѕ�t��   �M�ĝ����Pj�M��݊���ȅ�uW�}�u�U ����M ��@�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M�������P�M�U�}�u�E�   �w�}�t�}�u>�E�P�M$��Qjj�UR�EP�M�Q�+������U �M ��U$�B���M$�A�-�U�R�E$��Pjj�MQ�UR�E�P�������M �U ��EP�MQ赉�����Ѕ�t'�M�����PjH�M��ۉ���ȅ�t
�M�m����UR�EP�w������ȅ�t<j �M肜����R�M��eq���E��E��:t�M��,t	�U��/u�M�����EP�MQ�$������Ѕ�t'�M�1�����PjH�M��J����ȅ�t
�M�ܰ���UR�EP�]v�����ȅ�t�U ����M ��  �M������Rj�M����������uM�}�t�M ����E ��3�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��2�����P�M�U�   �}�u>�E�P�M$��Qjj�UR�EP�M�Q�X������U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P�������M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��2�����@�U�E�MQ�UR�u��������t�M ����E ��M�U��E�A�E�M�d�    Y��]�  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M�h}  h��EP�MQ�UR�EP谴����h~  h��M$Q�ٶ�����U��BPj �MQ�UR�X������E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U����M�h}  h��EP�MQ�UR�EP蚠����h~  h��M$Q�������U��BPj �MQ�UR膲�����E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M�h�   h��EP�MQ�UR�EP������h�   h��M$Q�:������U�R�M�ƍ���E�E�E��E�    �M�Q�ę�����E��E������M��f���U�R�E$��Pjj �MQ�UR�E�P�p�����M �U ��E �8 uj �M襂����Q�M��A����Ѓ�:t�E ����U �
�2�E�P�M$��Qj;j �UR�M�����P�E�P�$p�����M �U ��E �8 uj �M�>�����Q�M��ڄ���Ѓ�:t�E ����U �
�/�E�P�M$Qj;j �UR�M蛔��P�E�P��o�����M �U ��E�M��U�P�E�M�d�    Y��]�  ����������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P�����3�P�E�d�    �M�h�   h��EP�MQ�UR�EP苝����h�   h��M$Q�
������U�R�M薋���E�E�E��E�    �M�Q��f�����E��E������M��Xd���U�R�E$��Pjj �MQ�UR�E�P袕�����M �U ��E �8 uj �M脔����Q�M��gi���Ѓ�:t�E ����U �
�2�E�P�M$��Qj;j �UR�M����P�E�P�;������M �U ��E �8 uj �M������Q�M�� i���Ѓ�:t�E ����U �
�/�E�P�M$Qj;j �UR�M誨��P�E�P�ה�����M �U ��E�M��U�P�E�M�d�    Y��]�  ����������������������������������������������������������������������������������������������������������������������������U����M�hn  h��EP�MQ�UR�EP�Ю����ho  h��M$Q��������U��BPj �MQ�UR�x������E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U����M�hn  h��EP�MQ�UR�EP躚����ho  h��M$Q�9������U��BPj �MQ�UR覬�����E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U��j�h�d�    P�����3�P�E�d�    �M�h�  h��EP�MQ�UR�EP�1�����h�  h��M$Q�Z������U�R�M�����E�E�E��E�    �M�Q�������E��E������M��`���E�    �U�R�E�Ph�  j �MQ�UR�E�P�j�����M �U ��E ���u6�}�l  |�U���l  �U���}��   ~�E ����U �
�E$�M��H�U�E��M�J�E�M�d�    Y��]�  ��������������������������������������������������������������������������������U��j�hH�d�    P�����3�P�E�d�    �M�h�  h��EP�MQ�UR�EP�[�����h�  h��M$Q�ڭ�����U�R�M�f����E�E�E��E�    �M�Q��a�����E��E������M��(_���E�    �U�R�E�Ph�  j �MQ�UR�E�P�k������M �U ��E ���u6�}�l  |�U���l  �U���}��   ~�E ����U �
�E$�M��H�U�E��M�J�E�M�d�    Y��]�  ��������������������������������������������������������������������������������U����M��E�    �E��HQ�M�Σ���U����U��E��]� ���������������U����M��E�    �E��HQ�M莣���U����U��E��]� ���������������U����M��E�    �E��HQ�M�N����U����U��E��]� ���������������U����M��E�    �E��HQ�M�����U����U��E��]� ���������������U��Q�M�j{h���EP�MQ��������U+U����R�EP�R�������]� ���������������������U��Q�M�j{h���EP�MQ�9i�����U+U����R�EP��������]� ���������������������U����M�hq  h8��EP�MQ�`~����hr  h8��UR�EP��x�����M�U��E �M��U�;Eu	�E�    ��E�   �M��M�U�;E��   �M �;U��   �E��P�MQ�U�E+P�M�R�E �Q�W������E��U��U��}��t�}��t�}� t�4�E�M��E��]�   �V�U ����u�U�P�S��������E��}��u�E�    �M�U��E��M ����E ��E�    �8����E��]� ����������������������������������������������������������������������������������U����M�h�  h8��EP�MQ��|����h�  h8��UR�EP�7y�����M�U��E �M��U�;Eu	�E�    ��E�   �M��M�U�;E��   �M �;U��   �E��P�MQ�U�E+P�M�R�E �Q�ǫ�����E��U��U��}��t�}��t�}� t�4�E�M��E��]�   �V�U ����u�U�P�Ç�������E��}��u�E�    �M�U��E��M ����E ��E�    �8����E��]� ����������������������������������������������������������������������������������U��Q�M�hk  h8��EP�MQ������hl  h8��UR�������E���P�MQ�UR�EP�ds������]� ������������������������U����M��E���P�MQ�Ou�������E#�t	�E�   ��E�    �E���]� �������������������������������U��Q�M�h�
  h8��EP�MQ��d����h�
  h8��UR�������E���P�MQ�UR�EP�r������]� ������������������������U����M��E���P�MQ�t�������E#�t	�E�   ��E�    �E���]� �������������������������������U����M�h�  h8��EP�MQ�y�����U��E��E�    �M�M��U�;U��   �E�;E��   �M��Q�U�R�E+E�P�M�Q�U�R�֨�����E��E��E�}��t�}��t�}� t�$�E��F�E��A�M���u�U�R���������E��}��u�E�    �E�E��E��M���M��a����E��]� ����������������������������������������������������������������U����M�h�  h8��EP�MQ�x�����U��E��E�    �M�M��U�;U��   �E�;E��   �M��Q�U�R�E+E�P�M�Q�U�R趧�����E��E��E�}��t�}��t�}� t�$�E��F�E��A�M���u�U�R��������E��}��u�E�    �E�E��E��M���M��a����E��]� ����������������������������������������������������������������U��Q�M��   ��]�����������������U��Q�M��   ��]�����������������U��Q�M��EP�MQ�M���X����]� �����������������U��Q�M�h�  h8��EP�MQ��}����h�  h8��UR�U�������E���E�M���M�U;Ut�EP�M�R�M��OX���M��ˋE��]� �����������������������������������������U��Q�M��EP�MQ�M��Z����]� �����������������U��Q�M�h�
  h8��EP�MQ�`����h�
  h8��UR腓������E���E�M���M�U;Ut�EP�M�R�M��Y���M��ˋE��]� �����������������������������������������U��Q�M��E��H$�U�
�E��]� ���������������������U��Q�M��E��H$�U�
�E��]� ���������������������U����M��E�    �E��HQ�M�^���U����U��E��]� ���������������U����M��E�    �E��HQ�M�7y���U����U��E��]� ���������������U��Q�M������]� ����������������U��Q�M������]� ����������������U��� ���3ŉE��M�h�  h8��EP�MQ�1{����h�  h8��UR�EP�������M�U��E �M��U�;Eu	�E�    ��E�   �M�M�U�;E�  �M �;U�   蛘���M �U+;�]�E��P�MQ�U��Q�U �P�j������E��}� }�   �   �!�M����E��M �U��E ��E�    �   �M��U��E��P�MQ�U��Q�U�R�������E��}� }	�   �]�S�E �M+;M�}�U�E���E��A�7�M�Q�U�R�E �Q��]�����U����M��U �E��M ��E�    ������E�M�3��Is����]� ����������������������������������������������������������������������������������������������������������U��� ���3ŉE��M�h�  h8��EP�MQ��\����h�  h8��UR�EP�܏�����M�U��E �M��U�;Eu	�E�    ��E�   �M�M�U�;E�  �M �;U�   苖���M �U+;�]�E��P�MQ�U��Q�U �P�Z������E��}� }�   �   �!�M����E��M �U��E ��E�    �   �M��U��E��P�MQ�U��Q�U�R��������E��}� }	�   �]�S�E �M+;M�}�U�E���E��A�7�M�Q�U�R�E �Q��[�����U����M��U �E��M ��E�    ������E�M�3��9q����]� ����������������������������������������������������������������������������������������������������������U��Q�M��E��H �U�
�E��]� ���������������������U��Q�M��E��H �U�
�E��]� ���������������������U����M��E�    �E��HQ�M�aY���U����U��E��]� ���������������U����M��E�    �E��HQ�M��s���U����U��E��]� ���������������U��j�h��d�    P��d���3ŉE�P�E�d�    �M��E�P�M�{t���E��M��M��E�    �U�R�y������E��E������M��=M���E�P�   k�����R�   k� ����Q�M��:����E� �E�    �M ��~���Ѕ�u+j �M �6`��� �   k�
�L�;�u�E��U����U��M �����E��E��E��	�M����M��U�;U�s&�E�P�M ��_��f���R�E�P�՛������
s�ɋM�+M�Q�U�R�M �_��P�M������E�   �M��T~������t�   k� �D�Pj�M��"����   k� �D�P���̉e��U�R�{���E��E�P�MQ�UR�EP�MQ�UR�EP�M��e���E������M��u^���E�M�d�    Y�M�3��n����]� ����������������������������������������������������������������������������������������������������������������������������������U��j�h��d�    P��t���3ŉE�P�E�d�    �M��E� ���] ����Au�E��E ���] �E�    �	�E���
�E��E �(�����u�}��  s�E �5��] �Ѓ��E �$hH�j(�M�Q�W������E��}� }�U�E��M�J�E��   �U�R�M�q���E��E��E��E�    �M�Q�}�����E��E������M��MJ��j0�M��I]��f�E�j �U�R�M��6J���E�   j �M��	a��P�E��L�Q�   k� �L�Q�M��)����U�R�E�P�M��٘���M�Q���̉e��U�R��x���E��E�P�MQ�UR�EP�MQ�UR�EP�M��[c���E������M��5\���E�M�d�    Y�M�3���k����]�  ������������������������������������������������������������������������������������������������������������������U��j�h �d�    P��d���3ŉE�P�E�d�    �M��E�P�M��o���E��M��M��E�    �U�R�LK�����E��E������M��H���E�P�   k���P�R�   k� ��P�Q�M��~\���E� �E�    �M �O���Ѕ�u+j �M �L��� �   k�
�L�;�u�E��U����U��M 蝐���E��E��E��	�M����M��U�;U�s&�E�P�M �KL��f���R�E�P�m�������
s�ɋM�+M�Q�U�R�M �L��P�M���a���E�   �M��^N������t�   k� �D�Pj�M��N���   k� �D�P���̉e��U�R�U���E��E�P�MQ�UR�EP�MQ�UR�EP�M������E������M��dv���E�M�d�    Y�M�3��i����]� ����������������������������������������������������������������������������������������������������������������������������������U��j�hp�d�    P��t���3ŉE�P�E�d�    �M��E� ���] ����Au�E��E ���] �E�    �	�E���
�E��E �(�����u�}��  s�E �5��] �Ѓ��E �$hH�j(�M�Q�ǃ�����E��}� }�U�E��M�J�E��   �U�R�M��l���E��E��E��E�    �M�Q�\H�����E��E������M��E��j0�M��͔��f�E�j �U�R�M��R����E�   j �M���q��P�E��L�Q�   k� �L�Q�M��mY���U�R�E�P�M��iL���M�Q���̉e��U�R�eS���E��E�P�MQ�UR�EP�MQ�UR�EP�M��ތ���E������M��$t���E�M�d�    Y�M�3��Ag����]�  ������������������������������������������������������������������������������������������������������������������U���P���3ŉE��M��EP�M�ތ��Ph��M�Q�U�R��c����Pj@�E�P������P�M�Q�UR�EP�MQ�UR�EP�M�Q��U���� �E�M�3��Rf����]� �����������������������������������U���P���3ŉE��M��EP�M�>���Ph��M�Q�U�R�Oc����Pj@�E�P�O�����P�M�Q�UR�EP�MQ�UR�EP�M�Q�ZU���� �E�M�3��e����]� �����������������������������������U���   ���3ŉE���`����M茌����T�����X�����X��� 0|	��T��� w%�M�t���%    uǅh���   ǅl���    ��M�?�����h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M�����% 0  =    �  �E��^�E������D��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E�(�����u��x����  s�E�5��]���E�x^����Aud���t�����
��t����}� |M	��|���
rB���]����u2��t����  s&�E���]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M腉��Pj �E�P��`���Q�h����Pjl�U�R�~����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P�+�����,�E�M�3���b����]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE���`����M�,�����T�����X�����X��� 0|	��T��� w%�M����%    uǅh���   ǅl���    ��M�߈����h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M�`���% 0  =    ��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E�(�����u��x����  s�E�5��]���E�x^����Aud���t�����
��t����}� |M	��|���
rB���]����u2��t����  s&�E���]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M�>���PjL�E�P��`���Q�ee����Pjl�U�R�O{����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P������,�E�M�3��_����]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���H���3ŉE��M��EPh �j@�M�Q�)z����P�U�R�EP�MQ�UR�EP�MQ�U�R�4N���� �E�M�3��^����]� �����������������������������U���P���3ŉE��M��E P�MQ�M�z���Ph��U�R�E�P�[����Pj@�M�Q�y����P�U�R�EP�MQ�UR�EP�MQ�U�R�M���� �E�M�3���]����]� �����������������������������������������������U���P���3ŉE��M��E P�MQ�M�ʃ��Ph��U�R�E�P��Z����Pj@�M�Q��x����P�U�R�EP�MQ�UR�EP�MQ�U�R��L���� �E�M�3��>]����]� �����������������������������������������������U��j�h��d�    P��   ���3ŉE�VP�E�d�    �M�h�  h���EP��I�����M�����% @  u4�MQ�UR�EP�MQ�UR�EP�M���M��B$�ЋE��  ��  ��p���Q�M�;a���E��U���|����E�    ��|���P�g�����E��E�������p�����9���M��	����E�   �M��t%�U�R�M��A���E��E�P�M��es���M��ML���#�M�Q�M��UT���E��U�R�M��@s���M��(L���M�dg����t�����x�����x��� |:	��t��� v/�M�<g�����M�耇��;�v�M�&g�����M��j���+��u���E�    �E��E��M褁��%�  ��@t6�M�Q�UR�EP�MQ��`���R�E�P詈������P�M�U�E�    �M�����P�M��`��P�EP�MQ��h���R�E�P�Kf������P�M�Uj j �M�UL���E�P�MQ�UR�EP�MQ�U�R�2������E������M��K���E�M�d�    Y^�M�3��Z����]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������U���P���3ŉE��M��EP�M����Ph��M�Q�U�R�o����Pj@�E�P�u����P�M�Q�UR�EP�MQ�UR�EP�M�Q�y���� �E�M�3��Y����]� �����������������������������������U���P���3ŉE��M��EP�M�n��Ph��M�Q�U�R��n����Pj@�E�P�t����P�M�Q�UR�EP�MQ�UR�EP�M�Q�}x���� �E�M�3���X����]� �����������������������������������U���   ���3ŉE���`����M�����T�����X�����X��� 0|	��T��� w%�M�~��%    uǅh���   ǅl���    ��M�o����h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M��}��% 0  =    �  �E��^�E������D��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E�(�����u��x����  s�E�5��]���E�x^����Aud���t�����
��t����}� |M	��|���
rB���]����u2��t����  s&�E���]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M�|��Pj �E�P��`���Q��M����Pjl�U�R��q����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P�j����,�E�M�3��V����]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE���`����M�\|����T�����X�����X��� 0|	��T��� w%�M�D{��%    uǅh���   ǅl���    ��M�|����h�����l�����h�����|�����l����M��}� |	��|���$vǅ\���$   ���|�����\�����\�����p�����p������|���+ȋE��|����E�ǅx���    ǅt���    �M�z��% 0  =    ��   ���]����Auǅd���   �
ǅd���    ��d����M��U���t�E���]���x�����
��x����E�(�����u��x����  s�E�5��]���E�x^����Aud���t�����
��t����}� |M	��|���
rB���]����u2��t����  s&�E���]��|�����
�E��� ��|����E���M���t�E���]���E�$��p���R�M�ny��PjL�E�P��`���Q�J����Pjl�U�R�n����P��|���P��t���Q��x���R�E�P�MQ�UR�EP�MQ�UR��`���P�Wg����,�E�M�3���R����]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���H���3ŉE��M��EPh �j@�M�Q�Ym����P�U�R�EP�MQ�UR�EP�MQ�U�R�Wq���� �E�M�3��Q����]� �����������������������������U���P���3ŉE��M��E P�MQ�M�w��Ph��U�R�E�P� g����Pj@�M�Q�l����P�U�R�EP�MQ�UR�EP�MQ�U�R�p���� �E�M�3��Q����]� �����������������������������������������������U���P���3ŉE��M��E P�MQ�M��v��Ph��U�R�E�P�pf����Pj@�M�Q�l����P�U�R�EP�MQ�UR�EP�MQ�U�R�	p���� �E�M�3��nP����]� �����������������������������������������������U��j�h d�    P��   ���3ŉE�VP�E�d�    �M�h�  h���EP�y�����M� v��% @  u4�MQ�UR�EP�MQ�UR�EP�M���M��B$�ЋE��  ��  ��p���Q�M�kT���E��U���|����E�    ��|���P��-�����E��E�������p����$-���M��|^���E�   �M��t%�U�R�M���y���E��E�P�M���a���M���[���#�M�Q�M��R9���E��U�R�M���a���M���[���M�Z����t�����x�����x��� |:	��t��� v/�M�lZ�����M���t��;�v�M�VZ�����M���t��+��u���E�    �E��E��M��t��%�  ��@t6�M�Q�UR�EP�MQ��`���R�E�P�>l������P�M�U�E�    �M��xt��P�M��c��P�EP�MQ��h���R�E�P�W������P�M�Uj j �M�?���E�P�MQ�UR�EP�MQ�U�R��k�����E������M��Z���E�M�d�    Y^�M�3���M����]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h` d�    P��T���3ŉE�P�E�d�    �M�h&  h��EP�:����h'  h��MQ�X[�����L��U�P��E�f�T�f�M�M���[���E�    �U$��uf�E �   ��f�D��#f�U$�   ��f�T�f�M �   k�f�L��E�   ��M���M�j �U�R�M��1���M�����J��P�EP�M�Q�M��Nr��P�U�R�M��m���E��E��E��E��M��D7��P�if�����E��}� v	�E�   ��E�    �M��M��E� �M��?:���Uǅ�t��i����EP�MQ�U�R�M���U��Pj�M���U��P�EP�a�����E������M��YX���E�M�d�    Y�M�3��vK����]�  �����������������������������������������������������������������������������������������������������������������������U��j�h� d�    P��T���3ŉE�P�E�d�    �M�h�  h��EP�Ut����h�  h��MQ�(Y�����L��U�P��E�f�T�f�M�M��Y���E�    �U$��uf�E �   ��f�D��#f�U$�   ��f�T�f�M �   k�f�L��E�   ��M���M�j �U�R�M���.���M����H��P�EP�M�Q�M��p��P�U�R�M��uk���E��E��E��E��M��5��P�9d�����E��}� v	�E�   ��E�    �M��M��E� �M��8���Uǅ�t��i����EP�MQ�U�R�M��S��Pj�M��S��P�EP�<�����E������M��)V���E�M�d�    Y�M�3��FI����]�  �����������������������������������������������������������������������������������������������������������������������U��Q�M�ht  h8��EP�MQ�O�����	�U���U�E;Et�M�R�EP�M��o���ȅ�u�ҋE��]� ����������������������U��Q�M�h�
  h8��EP�MQ�V2�����	�U���U�E;Et�M�R�EP�M��\C���ȅ�u�ҋE��]� ����������������������U��Q�M�h}  h8��EP�MQ�=N�����	�U���U�E;Et�M�R�EP�M��/n���ȅ�t�ҋE��]� ����������������������U��Q�M�h�
  h8��EP�MQ�v1�����	�U���U�E;Et�M�R�EP�M��|B���ȅ�t�ҋE��]� ����������������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M��E�f�@��]���������������U��Q�M��E���P�MQ�=a������]� ���������������U��Q�M�h�  h8��EP�MQ�L�����	�U���U�E;Et�M���Q�U�P��`�����Mf��ыE��]� �������������������������������������U��Q�M�h�
  h8��EP�MQ��/�����	�U���U�E;Et�M���Q�U�P�^`�����Mf��ыE��]� �������������������������������������U��Q�M��E���P�MQ�`������]� ���������������U��Q�M��E���P�MQ�s������]� ���������������U��Q�M�h�  h8��EP�MQ�MK�����	�U���U�E;Et�M���Q�U�P�`s�����Mf��ыE��]� �������������������������������������U��Q�M�h�
  h8��EP�MQ�v.�����	�U���U�E;Et�M���Q�U�P��r�����Mf��ыE��]� �������������������������������������U��Q�M��E���P�MQ�r������]� ���������������U��j�hd�    P��\���3ŉE�VP�E�d�    �M��E�    jhh���EP�MQ��I�����M��Mr���E�    �U+U���Ũ}� ��   �E�P�M���b���M���Q�UR�EP�M�Q�M��)5���E��U��U��E��M��F�����M���n���FP�M�Q�M���4���E��U��U��E��M��VF��P�)�����E̍M��n��9E�w	�E�   ��E�    �EȈE��E��M��(���E� �M��(���MӅ�t��5����U�R�M��7b���E�P�M�� ���Mă��M��E������M��2���E�M�d�    Y^�M�3��QB����]� ��������������������������������������������������������������������������������������������������U��j�hXd�    P��\���3ŉE�VP�E�d�    �M��E�    jhh���EP�MQ�+�����M��P���E�    �U+U���Ũ}� ��   �E�P�M��zc���M���Q�UR�EP�M�Q�M���b���E��U��U��E��M��w,�����M��Ug���FP�M�Q�M��b���E��U��U��E��M��H,��P��m�����E̍M��g��9E�w	�E�   ��E�    �EȈE��E��M��</���E� �M��0/���MӅ�t��5����U�R�M��b���E�P�M�X���Mă��M��E������M��UM���E�M�d�    Y^�M�3��q@����]� ��������������������������������������������������������������������������������������������������U����M��E�    �E��HQ�M�)���U����U��E��]� ���������������U����M��E�    �E��HQ�M�C���U����U��E��]� ���������������U������3ŉE��M�h�  h8��EP�MQ�\�����U�E��E�    �M��U�E��P�MQj �U�R�sn�����E��}� 	�E�   �P�E����E��M�U+;U�}�E�M��E�   �)�}� ~#�U�R�E�P�M�R�T)�����E�M��U�
�E�M�3��>����]� ��������������������������������������������������������������U������3ŉE��M�h�  h8��EP�MQ�[�����U�E��E�    �M��U�E��P�MQj �U�R�cm�����E��}� 	�E�   �P�E����E��M�U+;U�}�E�M��E�   �)�}� ~#�U�R�E�P�M�R�D(�����E�M��U�
�E�M�3��=����]� ��������������������������������������������������������������U��Q�M��EP�M��8����]� ������U��Q�M�h�  h8��EP�MQ��<����h�  h8��UR��K������E���E�M���M�U;Ut�E�Q�M��K8���Uf��ϋE��]� �����������������������������U��Q�M�h�
  h8��EP�MQ�2<����h�
  h8��UR�=C������E���E�M���M�U;Ut�E�Q�M��T���Uf��ϋE��]� �����������������������������U��Q�M��EP�M��CT����]� ������U����M��E��x u	�E�   ��E�    �E���]������������������������U����M��E��x u	�E�   ��E�    �E���]������������������������U��Q�M��E�P�M��/���M��Q�PP�M��`���E��]� ������������������U��Q�M��E�P�M��HL���M��Q�PP�M�[���E��]� ������������������U����  ]�������U����  ]�������U��Q�E��U�;�u	�E�   ��E�    �E���]����������������������U��Q�E��U�;�u	�E�   ��E�    �E���]����������������������U����M��E��H��u�M�����U�B��u�M����M��9 u�U�: t�E��8 t�M�9 u	�E�    ��E�   �E���]� ����������������������������������������U����M��E��H��u�M���]���U�B��u�M�]���M��9 u�U�: t�E��8 t�M�9 u	�E�    ��E�   �E���]� ����������������������������������������U��Q�M��E��H;Ms�M��2���UR�M��>A���E���]� �����������������U����M��E��H;Ms�M��?2���U��B+E;Ew�MQ�M���@���L�} vF�M��-���U�P�E��M��Q+U�U�E�+EP�M�U��JP�M�Q�?�����U�R�M��@���E���]� �����������������������������������U��Q�M��E��H;Ms�M��6P���UR�M��	+���E���]� �����������������U����M��E��H;Ms�M���O���U��B+E;Ew�MQ�M��*���L�} vF�M���H���U�P�E��M��Q+U�U�E�+EP�M�U��JP�M�Q�"�����U�R�M��k*���E���]� �����������������������������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��E���M��B$�Ћ�]���������U��Q�M��E���M��B$�Ћ�]���������U����M��E�P�M��&��P�M�e���E��]� ���������U����M��E�P�M�����P�M��O���E��]� ���������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P �ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P �ҋE��]�  �������������������U��Q�M��E��H���]��������������U��Q�M��E��H���]��������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E��H;Ms�M��_,���U����+B;Ew�M��Q���} vx�M��QU�U�j �E�P�M�� ]���ȅ�tW�U��B+EP�M���&���M�HR�M���&���M�H�E�BQ�9�����UR�EP�MQ�M��,9���U�R�M��:���E���]� �����������������������������������������������������U����M��E��H;Ms�M��J���U��Ċ+B;Ew�M��|`���} vx�M��QU�U�j �E�P�M���%���ȅ�tW�U��B+EP�M���B���M�HR�M���B���M�H�E�BQ�������UR�EP�MQ�M��!���U�R�M��]$���E���]� �����������������������������������������������������U��Q�M��EP�MQ�U���M��P�ҋ�]� ������������U��Q�M��EP�MQ�U���M��P�ҋ�]� ������������U��Q�E���u	�E�    ��UR�;�����E��E���]��������������������U��Q�E���u	�E�    ��UR�t;�����E��E���]��������������������U��Q�M��E�P�D1������]����������U��Q�M��E�P�&������]����������U��Q�M�������]�����������������U��Q�M�������]�����������������U��M�8?��]����U��M��S��]����U����M��E�P�M��F��������E��}�w	�E�   �	�M����M�E��]�������������������U����M��E�P�M��������+H���E��}�w	�E�   �	�M����M�E��]�������������������U��Q�} u�E�E���MQ�UR�EP�W�����E��E���]�����������������U��Q�} u�E�E���MQ�UR�EP��V�����E��E���]�����������������U��j�h�d�    P��X���3ŉE�P�E�d�    �M��E�    �E��8 u)�M��wZ���E��M��M��E�    �U����U��E��E��(�M��	����>��P�M��Q���E��U����U��E��E��M��M��U�R�M�����E����E��M���t�e���M��#���E������U���t�e���M�����E�M�d�    Y�M�3��-����]� �������������������������������������������������������������U��Q�M��EP�MQ�U���M��P8�ҋ�]� ������������U��Q�M��EP�MQ�U���M��P8�ҋ�]� ������������U��Q�M��EP�M���M��B,�ЋE��]� ���������������U��Q�M��EP�M���M��B,�ЋE��]� ���������������U����M��E�    �EP�M���M��B �ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B �ЋM����M��E��]� �������������U��Q�M��EP�M���M��B(�ЋE��]� ���������������U��Q�M��EP�M���M��B(�ЋE��]� ���������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E��H;Mr�M�W��;Es�M��$���U��B+E;Es�M��Q+U�U�M��V��+E�E��E�;Es�M��M���+U�E��H+M;�w�M��I���U��B+E+E�E��M��QU+U�U�E��H;M�sj �U�R�M���T���E�;Ete�M�Q�M������U�P�M�HR�M������M�H�E�BQ�1�����UR�M�t���M�HR�M�����M�HR�������  �E;Ewe�MQ�M��j���U�PP�M��[���M�HR�(1�����E�P�M��@���M�H�E�BQ�M��+���U�P�M�HR��0�����|  �E;Ewe�M�Q�M������U�P�M�HR�M������M�H�E�BQ�0�����UR�M������M�HR�M�����M�HR�0�����  �EE;Ewk�M�Q�M�����U�P�M�HR�M��x���M�H�E�BQ�?0�����UR�M��W���MM+M�HR�M��B���M�HR�0�����   �EP�M��"���M�HR�M�����M�HR��/�����E�P�M������M�H�E�BQ�M������U�P�M�HR�/�����E+EP�M�����M�H�E�BQ�M�����U�P�M�HR�q/�����E�P�M��a0���E���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��} th�  hXo�EP�N/�����MQ�M��zN���Ѕ�t-�EP�M��h���M+���Q�U�R�EP�MQ�M�����5  �U��B;Es�M��C ���M��Q+U;Us�E��H+M�M���+U�E��H+M;�w�M���D���U��B+E+E�E��M;Ms6�U�R�M������M�H�E�BQ�M������U�P�M�HR�-�����} w
�} ��   �E��HM+M�M�j �U�R�M��mP������ti�M;Ms6�U�R�M��j���M�H�E�BQ�M��U���U�P�M�HR�-�����EP�MQ�M��0���U�PP�\�����M�Q�M���-���E���]� ����������������������������������������������������������������������������������������������������������������U��j�h9d�    P��   ���3�P�E�d�    �M��E�   �E,P�M �,���ȅ���   ���̉e��UR��R���EȋEȉE��E����̉e��UR��R���E��E��+�����EЋE�P��p���Q�M�����E��U��U��E����̉e��E�P�R���E؋M؉M��E����̉e��UR�zR���E��E��E+�����E�E�P�M��U���E���p����Y
����   �M Q�M,�A%��P�M �'��P���̉�|����UR�R���E�E�E��E����̉e��UR� R���E��E���*�����E�E�P��d���Q�M������E܋U܉U��E����̉e��E�P�Q���E̋M̉M��E�	���̉e��UR�Q���E��E��j*�����EċE�P�M��2���E���d����~	���M��M��E��M�	���E��M�	���E� �M �T	���E������M,�E	���E��M�d�    Y��]�0 ��������������������������������������������������������������������������������������������������������������������������������������������������U����M��E��H;Mr�M�H��;Es�M��g:���U��B+E;Es�M��Q+U�U�M�nH��+E�E��E�;Es�M��M���+U�E��H+M;�w�M��P���U��B+E+E�E��M��QU+U�U�E��H;M�sj �U�R�M������E�;Ete�M�Q�M���2���U�P�M�HR�M���2���M�H�E�BQ�������UR�M�G2���M�HR�M��2���M�HR��������  �E;Ewe�MQ�M��y2���U�PP�M��j2���M�HR�a�����E�P�M��O2���M�H�E�BQ�M��:2���U�P�M�HR�+�����|  �E;Ewe�M�Q�M��2���U�P�M�HR�M���1���M�H�E�BQ�������UR�M���1���M�HR�M���1���M�HR������  �EE;Ewk�M�Q�M��1���U�P�M�HR�M��1���M�H�E�BQ�x�����UR�M��f1���MM+M�HR�M��Q1���M�HR�H�����   �EP�M��11���M�HR�M��"1���M�HR������E�P�M��1���M�H�E�BQ�M���0���U�P�M�HR��
�����E+EP�M���0���M�H�E�BQ�M��0���U�P�M�HR�
�����E�P�M��\���E���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��} th�  hXo�EP��#�����MQ�M�����Ѕ�t-�EP�M��w/���M+���Q�U�R�EP�MQ�M��J���5  �U��B;Es�M��(6���M��Q+U;Us�E��H+M�M���+U�E��H+M;�w�M��sL���U��B+E+E�E��M;Ms6�U�R�M���.���M�H�E�BQ�M���.���U�P�M�HR�������} w
�} ��   �E��HM+M�M�j �U�R�M��f������ti�M;Ms6�U�R�M��y.���M�H�E�BQ�M��d.���U�P�M�HR�U�����EP�MQ�M��?.���U�PP������M�Q�M������E���]� ����������������������������������������������������������������������������������������������������������������U��j�h�d�    P��   ���3�P�E�d�    �M��E�   �E,P�M � H���ȅ���   ���̉e��UR�S���EȋEȉE��E����̉e��UR�5���E��E��o�����EЋE�P��p���Q�M��=���E��U��U��E����̉e��E�P�����E؋M؉M��E����̉e��UR�����E��E�������E�E�P�M�������E���p�����	����   �M Q�M,�7��P�M ���P���̉�|����UR�x���E�E�E��E����̉e��UR�Z���E��E�������E�E�P��d���Q�M��<���E܋U܉U��E����̉e��E�P����E̋M̉M��E�	���̉e��UR�����E��E��3�����EċE�P�M�����E���d����	���M��M��E��M�u����E��M�i����E� �M �����E������M,�����E��M�d�    Y��]�0 ��������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M�j �EP�M��g!����]� ���������������������U��Q�M��E��M;Hw�UR�M��!����EP�M��U+QR�M��F����]� �������������������U��Q�M�j �EP�M��7����]� ���������������������U��Q�M��E��M;Hw�UR�M�������EP�M��U+QR�M�������]� �������������������U����M��M���%���E��U�}� |�}� v�M������P������f�E���E���M��B��f�E�f�E���]����������������������������U����M��M���B���E��U�}� |�}� v�M���>��P������f�E���E���M��B��f�E�f�E���]����������������������������U����M��E�P�M�Q�B����P�M�R���E��]� ���������������������U����M��E�P�M�Q��G����P�M�6���E��]� ���������������������U��Q�M��E�P�M��E���E��]� ��������������������U��Q�M��E�P�M�0���E��]� ��������������������U��EP�M������E]�������������U��EP�M�A���E]�������������U����M��M���#���E��U�}� |�}� v�M�� ��P������f�E���E���M��B��f�E�f�E���]����������������������������U����M��M���@���E��U�}� |�}� v�M��)B��P������f�E���E���M��B��f�E�f�E���]����������������������������U��Q�M��E��@��]����������������U��Q�M��E��@��]����������������U����M��M��s@���E�U��}� |/�}� v'�M������E�E�f�Mf��U�R�����f�E��!�EP�������Q�U���M��P��f�E�f�E���]� �����������������������������������������U����M��M�����E�U��}� |/�}� v'�M�� ���E�E�f�Mf��U�R�z����f�E��!�EP�h������Q�U���M��P��f�E�f�E���]� �����������������������������������������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Ef� ]������U��Ef� ]������U��Ef� ]������U��Ef� ]������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��EP�M���M��B0�Ћ�]� �����������������U��Q�M��EP�MQ�UR�E���M��B,�Ћ�]� ����������U��Q�M��EP�MQ�UR�E���M��B,�Ћ�]� ����������U��Q�M��EP�M���M��B0�Ћ�]� �����������������U��E��P�MQ�UR�������]����������������������U��E��P�MQ�UR�������]����������������������U��Q�E�E���M����M��U���U�} v�E�f�Mf��܋E��]��������������������������U��Q�EP�MQ�	�����E��U�R�EP�MQ�UR�EP�MQ�������E��]������������������U��Q�EP�M�Q�/������UR�E�P������M�Q�U�R�EP�MQ�UR�EP�MQ�L������E��]��������������������������������U����M�y����E���E�M;Mt�U�P�M�9������@���ϋM�U��E�A�E]������������������������U��EP�MQ�UR�EP�MQ�������E]�������������U����M��E��H(��t�U�B�E��	�M�Q�U��E���,Pj �M�Q�V������U��B�E�H.��v	�E��Q�	�U�B �E�M���,Qj �U�R�������M��A�U�B/��v	�E��	�M�Q$�U��E���,Pj �M�Q��������U��B�E���,Pj �   k� �E�H�R�.������M��A�U���,Rj �   k� �U�B�Q�������U��B��]� ���������������������������������������������������������������������������������U���4���3ŉE�VW�M̍E�P�M�C#���}̃��   ���M̃�Qj �M����P��������ỦB�Ẽ�Pj �M�����P��������M̉A�Ũ�Rj h���������M̉A_^�M�3������]� ��������������������������������������������������U��Q3��E��E���]�����������������U��E]���������U��EP�MQ�UR�EP�MQ�3����]����������������U��EP�MQ�UR�EP�MQ�=9����]����������������U��Q�E���]������U��E]���������U��j�hXd�    P��`���3�P�E�d�    �M��E�   ���̉eȍEP�����E�M�M��E����̉e��UR����E�E�E��E��M�Q�M������E�U�U��E����̉e��E�P�����E܋M܉M��E��U�R�M�����E؋E؉E��E����̉e��U�R����E��E��M��u(���EЋEЉE��E��M��	���E��M��	���E� �M�	���E������M�	���E̋M�d�    Y��]� �������������������������������������������������������������������������������������U��Q�E;Eu�M�U��E�A�E�{�yhQ  h8��MQ�UR�()����hR  h8��EP� �����MQ�UR������E��E�P�MQ�UR�EP������P�MQ�����P�UR�������E��]���������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M������E�    �P��E�0������E�M�Q�M�	���E�}� t�n�}� t�U��U��`�EP�M�Q���������uh|]�M�����hH=�U�R�����.�E��E�M��P��U��U�E��M�B�ЋM�Q�{)�����U�U��E������M��7#���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M��[����E�    �T��E�4��x����E�M�Q�M�����E�}� t�n�}� t�U��U��`�EP�M�Q�"��������uh|]�M��k���hH=�U�R����.�E��E�M��T��U��U�E��M�B�ЋM�Q�;(�����U�U��E������M���!���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M������E�    �X��E�8��8����E�M�Q�M����E�}� t�n�}� t�U��U��`�EP�M�Q�4��������uh|]�M��+���hH=�U�R�o���.�E��E�M��X��U��U�E��M�B�ЋM�Q��&�����U�U��E������M�� ���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h(d�    P��$���3�P�E�d�    j �M�������E�    �\��E�<�������E�M�Q�M�I���E�}� t�n�}� t�U��U��`�EP�M�Q�T(�������uh|]�M������hH=�U�R�/���.�E��E�M��\��U��U�E��M�B�ЋM�Q�%�����U�U��E������M��w���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�hXd�    P��$���3�P�E�d�    j �M������E�    �d��E�D������E�M�Q�M�	���E�}� t�n�}� t�U��U��`�EP�M�Q��������uh|]�M�����hH=�U�R�����.�E��E�M��d��U��U�E��M�B�ЋM�Q�{$�����U�U��E������M��7���E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M��[����E�    �`��E�@��x����E�M�Q�M�����E�}� t�n�}� t�U��U��`�EP�M�Q�J(�������uh|]�M��k���hH=�U�R����.�E��E�M��`��U��U�E��M�B�ЋM�Q�;#�����U�U��E������M������E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M������E�    �h��E�H��8����E�M�Q�M����E�}� t�n�}� t�U��U��`�EP�M�Q����������uh|]�M��+���hH=�U�R�o���.�E��E�M��h��U��U�E��M�B�ЋM�Q��!�����U�U��E������M�����E܋M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    j �M�������E�    �l��E�L�������E�M�Q�M�I���E�}� t�n�}� t�U��U��`�EP�M�Q�#�������uh|]�M������hH=�U�R�/���.�E��E�M��l��U��U�E��M�B�ЋM�Q� �����U�U��E������M��w���E܋M�d�    Y��]��������������������������������������������������������������������������U��Q�M��EP�M�����E���]� ��������������������U��j�hd�    PQ���3�P�E�d�    �M��EP�M��)���E�    �M��l��U��E�B(�MQ�UR�M��� ���E������E��M�d�    Y��]� �����������������������������������������U��Q�M��EP�M��K����M��U�B�A�E���]� ������������������������U��Q�M��M�����E��@    �E���]�����������������U��Q�M��EP�M�����E���]� ��������������������U��j�hHd�    P�����3�P�E�d�    �M�M��&��P�M�������E�    j j �M�� ����EP�MQ�M������E������E�M�d�    Y��]� �����������������������������������������U��j�hxd�    PQ���3�P�E�d�    �M��EP�M��<����E�    �M�����UR�M��t/���E������E��M�d�    Y��]� ���������������������������������������U��j�h�d�    PQ���3�P�E�d�    �M��EP�M��$���E�    �M����UR�M��N.���E������E��M�d�    Y��]� ���������������������������������������U��j�h�d�    PQ���3�P�E�d�    �M��EP�M������E�    �M��4��UR�M��L���E������E��M�d�    Y��]� ���������������������������������������U��j�hd�    PQ���3�P�E�d�    �M��EP�M������E�    �M��P��UR�M��k����E������E��M�d�    Y��]� ���������������������������������������U��Q�M��EPj�MQ�UR�M��_����E�� ��E���]� ����������������U��Q�M��EPj �MQ�UR�M������E�� ���E���]� ����������������U��j�h8d�    PQ���3�P�E�d�    �M��EP�M��6����E�    �M��,��UR�M������E������E��M�d�    Y��]� ���������������������������������������U��j�hsd�    PQ���3�P�E�d�    �M��EP�M�������E�    �M��`�j �M��������E��UR�M������E������E��M�d�    Y��]� ��������������������������������������U��Q�M��E�� l��M���%���M�������]�������������U��Q�M��E�� ���M��QR�T!�����M�������]����������������������U��Q�M��E�� ��M��	����]���������������������U��Q�M��E�� 4��M��R�����]���������������������U��Q�M��E�� P��M��"�����]���������������������U��Q�M��E�� ��M��
����]���������������������U��Q�M��E�� ���M��d
����]���������������������U��Q�M��E�� ,��M��*���M��l����]�������������U��Q�M��E�� `��M����"���M��W�����]����������U��Q�M��EP�M������E���]� ��������������������U��Q�M��EP�M������M��U�B�A�E���]� ������������������������U����M��E�;E��   j j�M��k���3�t�U�R�M���P�M������E�P�M���P�M�Q�M�����P��������Ѕ�t,���ĉe�P�M�?������̉e�Q�M�Z
���M�������UR�f����P�M������E���]� ���������������������������������������������������U����M��EP�M��5����M��U�A;Bu	�E�   ��E�    �E���]� ��������������������U����M��EP�M��&���ȅ�u	�E�   ��E�    �E���]� ���������������������������U��QV�M��M��������t-�E��x t$�M����������������M�����p�M�;qw_jmhXohH��O������ Y��t3�u#hPYh�Yj jnhXoj�P�������u�j jnhXoh��h�Z�������U��B���M��A�E�^��]����������������������������������������������������������U��Q�M��E���]� ����������������U��Q�M��EP�M������M��U�A+B��]� �����������U��j�h�d�    P�����3�P�E�d�    �M��E�    �E�P�M������E�    �MQ�M�����P�M�r����U����U��E������M�������E�M�d�    Y��]� ���������������������������������������������U��j�h�d�    P�����3�P�E�d�    �M��EP�M�Q�M��-���E�U�U��E�    �M������E��E������M��j����E�M�d�    Y��]� ������������������������������������������U��j�hd�    P�����3�P�E�d�    �M��E�    �E�P�M��>����E�    �MQ�M��n��P�M�"����U����U��E������M������E�M�d�    Y��]� ���������������������������������������������U��QV�M��M�������tN�E��x tE�M��qu�M��{���������;�r)�M��h������������M��W���p�U��BE;�shh�   hXohH��������� Y��t3�u&hPYh�Yj h�   hXoj���������u�j h�   hXoh��h�Z������M��QU�E��P�E�^��]� �������������������������������������������������������������U��Q�M��EP�M��1���E���]� ��������������������U��Q�M��E��P�M������]� ���������������������U��Q�M��M��-���E��t�M�Q�A������E���]� ��������������������U��Q�M��M�������E��t�M�Q�������E���]� ��������������������U��Q�M��M��v����E��t�M�Q��������E���]� ��������������������U��Q�M��M��o����E��t�M�Q�������E���]� ��������������������U��Q�M��M������E��t�M�Q�A������E���]� ��������������������U��Q�M��M������E��t�M�Q�������E���]� ��������������������U��Q�M��M��e!���E��t�M�Q��������E���]� ��������������������U��Q�M��M�����E��t�M�Q�������E���]� ��������������������U��Q�M��M��K���E��t�M�Q�A������E���]� ��������������������U��QV�M��M��������t�M���������M�����;�thh�   hXoh���c���������t3�u&h�h�Yj h�   hXoj�a�������u�j h�   hXoh��hx������^��]� ���������������������������������������U��j�h}d�    P��x���3ŉE�P�E�d�    �E�    �} ��   �E�8 ��   ����E�jChX��M�Qj�������E��E�    �}� tbj �U�R�M������E��E��E��E��MЃ��MЋM��\���P��|����p����E��U��U��E�   �EЃ��EЋM�Q�M�����E���E�    �UȉU��E�   �E�M���E�   �UЃ�t�e����|�������E������EЃ�t�e���M�������   �M�d�    Y�M�3�������]������������������������������������������������������������������������������������������U��j�h�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �x���E�jMh��M�Qj��������E��E�    �}� t:j �M�b��P�M�������E��U��U��E��E����E��M�Q�M�������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]�����������������������������������������������������������������������������U��j�hTd�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �8���E�h�  h��M�Qj�������E��E�    �}� t:j �M���P�M������E��U��U��E��E����E��M�Q�M��j����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h�d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �� ���E�h�  h��M�Qj�_������E��E�    �}� t:j �M����P�M��u����E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]��������������������������������������������������������������������������U��j�h4	d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �����E�h(  h��M�QjX�������E��E�    �}� t<jj �M���P�M��3����E��U��U��E��E����E��M�Q�M��|����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M��K���   �M�d�    Y��]������������������������������������������������������������������������U��j�h�	d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �x����E�h(  h��M�QjX��������E��E�    �}� t<jj �M�] ��P�M�������E��U��U��E��E����E��M�Q�M��L����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]������������������������������������������������������������������������U��j�h
d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   �8����E�h�   h���M�QjD�������E��E�    �}� t:j �M����P�M������E��U��U��E��E����E��M�Q�M��#����E���E�    �U�U��E�   �E�M؉�E������U���t�e���M������   �M�d�    Y��]��������������������������������������������������������������������������U��j�h�
d�    P��P���3�P�E�d�    �E�    �} ��   �E�8 ��   ������E�h�  h���M�Qj�_������E��E�    �}� t:j �M�����P�M��u����E��U��U��E��E����E��M�Q�M������E���E�    �U�U��E�   �E�M؉�E������U���t�e���M�����   �M�d�    Y��]��������������������������������������������������������������������������U��j�h�
d�    P�����3�P�E�d�    �M��E�P�M�����E�M�M��E�    �U�R�������E��E������M�������	�E(���E(�M(�����   �E(���%uO�U(���U(j �E(�Q�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M���M��B$�Ћ�P�M�U�   �E(��� uB��M������UR�EP��������ȅ�t�M�F�����RjH�M��q�������t���<j �M�#�����Q�M�������ЋE(�;�t�U ����M ����M�t��������UR�EP�;������ȅ�t�U ����M ��U�E��M�J�E�M�d�    Y��]�$ �����������������������������������������������������������������������������������������������������������������������U���@���3ŉE��E܉EԋMQ�UR�h���������t�[j �M�������Q�M �����E��Uۃ�+u�E�� +�Mԃ��MԋM�J���� �Uۃ�-u�E�� -�Mԃ��MԋM�(����E� �UR�EP�������ȅ�t,j �M������R�M �'�������0u�E��M�������Mڅ�t�U��0�Eԃ��EԹ   k��D܉E���E��M�����MQ�UR����������tFj �M�	�����Q�M �����E��Uۃ�0|$�Eۃ�9�MԊUۈ�E�;E�s	�Mԃ��M���Uڅ�u�E܉EԋM�� �E�    �U�Rj
�E�P�M�Q�u������E��E�    �UR�EP��������ȅ�t	�UЃ��UЍE�9E�t�}� u�M�;M|�U;U�}�EЃ��E���M�Ủ�EЋM�3��^�����]����������������������������������������������������������������������������������������������������������������������������������U��j�hJd�    P��  ���3ŉE�VP�E�d�    ������ǅ|���    h�  h(��E�HQ�R�E�HQ�R��
�����E��tQ������Q�M�)���������������������E�    �����P���������p����E������������ٽ���O������Q�M������������������������E�   ������P��������p����E�����������舽��ƅ���� ƅw��� �M������E�   ��D���Q��p��������M�����E�������R�M�N����������������������E�������Q���������4����E������������UR�   k�����Q�   k� ��P��4����
���ǅX���    ���X�������X������������D  ��X����7  ��X�����D�����L�����L����� ��L�����L���X�  ��L�����s�$��r�U�R��p����Z����E�������D����E��M�����u=�EP�MQ�������Ѕ�t&�M�,������M��l���� ;�tj �M�������Q��X���uH�M��4�����w;�MQ�UR�G���������u�M��������M������;�t
j �M�������x���R�M������������������������E�������Q�����������E���x�������������������M������UR�EP��������ȅ�tv��l���R�M�� ��������������������E���|�������|���������R��������������t)�M������������������;�uǅ8���   �
ǅ8���    ��8�����_����E�   ��|�����t��|������l����������_�����t������T���R�M��@����������������������E�	������Q������L�����T����E���T����{�����T�����tƅ�����E�������k����E��M��p����  �EP�MQ�\������Ѕ�t�t  ������P��p��������������������� ����E�
��|�������|����� ����������vej ������P��p����p����������������������E�   ��|�������|����������i����0�M�Y�����;�uǅ$���   �
ǅ$���    ��$�����g����E�
   ��|�����t��|�����������j����E�   ��|�����t��|�����������F�����g�����t?�M�X���������R��p�������������������P�M�����������������!  ��,���Q��p����0����������������������E���|�������|���������������vej �����Q��p��������������������������E�   ��|�������|��������������0�M������;�uǅ(���   �
ǅ(���    ��(�����f����E�   ��|�����t��|�����������E�   ��|�����t��|������,����������f�����tF�M����������P��p�������������������Q�M��m�������������ƅw�����   ������R��p��������������������X�����uǅ0���   �
ǅ0���    ��0�����U����������N�����U�����t�f��H���R��p����u����������������������uǅ<���   �
ǅ<���    ��<�����W�����H����������W�����tƅw�����  ǅ`���    ��p����������H�����d���R��p���������E���d����s�����u	ƅo��� ���p����������o�����o�����n�����n�����t��d����G������|e��M�m����EP�MQ�^������Ѕ�t?�M�������P�MQ���������h�����h���
s��h�������P�M�������L  j j�M��s����E�ǅx���    ��M�����MQ�UR�������������   �M�H�����Q�UR�y�������h�����h���
sV��h�������Q�M�������x���R�M��	���� ��t'��x���Q�M�������,�����,������,�����K��x���R�M��ɿ��� ��t�M��������n���;�t�"�j j�M��������x�������x���������x��� u�.��x���Q�M��n������~��x�������x����ƅ������d���芿����P�������������   ��x��� ��   ��P������u
�   �   ��x�������x���t��P����2��x���P�M������;�u(��x��� u(��P����2��x���P�M�蹾���;�}	ƅ�����%�   �� ��P������~��P�������P����A�����������t �E��M�������E���d���������  �E��M�������p����D�����l����MQ�UR������������   ��l�������   �M� �������l���;���   �MQ�M�e���P�]������Ѕ�t\��`���;�H���}N�M������Q�UR���������h�����h���
s'��h�������Q�M�������`�������`���눋�`���;�H���}ƅ�����M�������u	ƅ�����+���`�������`�����`���;�H���}j0�M�誽�����E���d����p����   ��X���u�vƅm��� ��M�t����EP�MQ�e������Ѕ�t)�M�������PjH��4���������ȅ�t	ƅm���븋�X�����D����� u��m�����uƅ������������������  �M���������  ������D����E���<���P�M��9����������������������E�������R����������E���<����N�����M苻����`���P�M������������������������E���|����� ��|���������P������3�����賹���ȅ�t@�UR�EP�(������ȅ�t)�M����������������;�uǅ@���   �
ǅ@���    ��@�����e����E�   ��|����� t��|���ߍ�`����v�����e�����t������H���P�M��߿���������������������E�������R�����������V����E���H���������V�����tƅ�����E�������
�����������tj �M��������w�����tj-jj �M������E�P�M�v�����|�����@��|����E��M�������E������M������E�M�d�    Y^�M�3��h�����]� �"p�e"h�k�p  �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��E�    �6���P�M�8����E����E��E��]� ����������������U��j�h�d�    PQ��@���3ŉE�SVWP�E�d�    �e��M��E�P�M������}���,�   ���M�����E��M��A    �U��B    �E��@    �M��A    �E�    �U���,Rj �E��HQ�4������E��U��E��B�M�Qj �M��J�����M�����j j �3����{x��E�������E������U��B(��t�M��Q(�U��	�E��H)�M��U��E��P�M��y |	�U��z|
�E��@    �M��Q.R�E��H*Q�U��B+P�M��� Q�M��7����U��B/P�M��Q,R�E��H-Q�U���$R�M������E��t,jh ��M��� Q裵����jh ��U���$R荵�����M�d�    Y_^[�M�3��������]� �������������������������������������������������������������������������������������������������������������������������U����M��E�P�M������P�E��H�P��]� �����������������������U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��j�hd�    PQ��SVW���3�P�E�d�    �e��M�E��@    �M��A    �U��B    �E�    �EPj �M��L����M�����E�M�U�Q��M��]���j j �������z��E�������E������M�d�    Y_^[��]� ���������������������������������������������U��j�hHd�    P�����3�P�E�d�    �M�E�P�M�7����E��M��M��E�    �U�R�M��� ����E������M��5����M�d�    Y��]� �����������������������������U��j�h3d�    P��   ���3�P�E�d�    j j �j������   ������#Uu�   �} um������E�j'h؝�E�Pj�5������E��E�    �}� tj �MQ�M������E���E�    �U�U��E������0�裱��P�E�P�M����� �0�花��P�MQ������P�M�y���j j �J������   ������#Uu�   �} um�����E�j(h؝�E�Pj聸�����E��E�   �}� tj �MQ�M������E���E�    �U�U��E������4�����P�E�P�M����� �4��ְ��P�MQ�=�����P�M�ſ��j j �������   ������#Uu�   �} um�c����E�j)h؝�E�Pj�ͷ�����E��E�   �}� tj �MQ�M�迮���E���E�    �U܉U��E������8��;���P�E�P�M�3���� �8��"���P�MQ轰����P�M����j j �������   ������#Uu�   �} um�����E�j*h؝�E�Pj�������E��E�   �}� tj �MQ�M�������E���E�    �UԉU��E������<�臯��P�E�P�M����� �<��n���P�MQ������P�M�]���j j �V������   ������#Uu�   �} uo������E�j+h؝�E�PjX�e������E��E�   �}� tj j �MQ�M�������E���E�    �ỦU��E������@��Ѯ��P�E�P�M�ɽ��� �@�踮��P�MQ������P�M觽��j j �$������   ������#Uu�   �} uo�E����E�j,h؝�E�PjX诵�����E��E�   �}� tj j �MQ�M��3����E���E�    �UĉU��E������D�����P�E�P�M����� �D�����P�MQ�������P�M����j j �������   ������#Uu�   �} us�����E�j-h؝�E�PjD��������E��E�   �}� tj �MQ�M�褬���E���E�    �U���|����E������H��d���P��|���P�M�Y���� �H��H���P�MQ������P�M�7���j j �j������   ������#Uu�   �} uy�������x���j.h؝��x���Pj�9������E��E�   �}� tj �MQ�M�������E���E�    �U���t����E������L�褬��P��t���P�M虻��� �L�般��P�MQ�Z�����P�M�w����M�d�    Y��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��E��H(��u,�}w&�}w �}wkU�E��kU(�����E���E� ��M��M�j�U�Rj�EP���������]� �������������������������U��j�h�d�    P�����3�P�E�d�    �E�   �} u	�E�    ��EP�M�����E��M��M��E� �M�p����E������M�a����E�M�d�    Y��]������������������������������������U��j�h�d�    P���3�P�E�d�    �E�    ��E ���E �M�J����M�����}  v�M�������R�M�S�����������E�M��U�P�E������M覦���E�M�d�    Y��]�����������������������������������������U��j�h�d�    P��  ���3ŉE�P�E�d�    ��X����E�    h  h(��EP�������M��tK������R�M�����������������������E�������Q�h�������8����E� �������c����I��t���R�M�b�����������������|����E���|���Q�:�������8����E� ��t��������U�R��8���������E���8����z������������� }������؉����������������������@����M$����;�@���w(�E@P�M$�������@���+ȃ�Qj �M$�3�����   �M����������   �M��צ��� ����   ��8����$�����/����M�賦����0����M$葰��+�@�����(�����0������tx��0������~k��0����;�(���sZ��0������(���+�(�����/���Qj��(���R�M$�x����   �� ��0������~��0�������0����z����M�������E��M ��tH��`���R��8����:���� ������M�Q��8����/�����x�����x���R�M������M��̫���L��H���P��8���������������H���R��8�������������������P�M��=�����H����~����M��R����E��M�j�����t2��d���Q��8�������������������R�M��������d����3���ƅ?��� ǅD���    ǅ4���    ���4�������4�����4����  ��4����������$�����$����� ��$�����$���X��   ��$�������$����M�臮���D�����D����   �M��n����D�����D����   ��@��� vǅ���   �
ǅ���    �M$�6���;�@���w�M$�&�����@���+ȃ�������
ǅ���    �M$�������������D�����D������D�������D�����4���tƅ?���������M�>��������������������� |1	������ v&�M����;�D���v�M����+�D���������
ǅ���    �������D����M�~���%�  ����������@tO�����   u��?�����u8��D���R�EP�MQ�UR������P�*�������P�M�UǅD���    ǅ4���    ���4�������4�����4����  ��4���������� ����� ����� �� ����� ���X��  �� ��������$�l��M�耬��P�����P�M��)����������������������E����̉�@���������R�������8����EP�MQ������R��������������������P�M�U�E�����������5  �M���������   j��$���P�M������������������������E����̉�0���������R�\�����L����EP�MQ������R��������������������P�M�U�E���$����o����  ��@��� ��   �M$�P���P�����P�M$������������������������E����̉�P���������R�������p����EP�MQ������R���������������������P�M�U�E�������մ���  �M$�ê��;�@����	  �E@Pj �M�������>�����������8����d�����Qj �M�\����������������M$�k�����@���+�R�E@P�MQ�UR��|���P�g�������P�M�U�M$�3���P������P�M$������������������������E�	���̉�d���������R������<����EP�MQ��l���R���������������������P�M�U�E�������踳���y  �M$覩��+�@���P������P�M$�I����������������������E�
���̉�\���������R������D����EP�MQ��t���R�6�������������������P�M�U�E��������%�����8���������Pj �M�������������������@���Q��@���R������P������Q�M$�b����������������������E�������������������������������E����̉�T���������R�6�����4����EP�MQ������R�Z�������������������P�M�U�E��������I����E��������:����mj�EP�MQ�UR������P�6�������P�M�U�����   u8��D���P�MQ�UR�EP������Q���������@�U�EǅD���    ������M�蹧������   �M�訧����Pj�� ���Q������R�M��E����������������� ����E��� ���������������������������E����̉�l���������R�������h����EP�MQ������R��������������������P�M�U�E��� ���� ����E�����������j j �M�<�����D���P�MQ�UR�EP�MQ�������E��M��ۢ���E��M��Ϣ���E� �M��â���E������M$财���E�M�d�    Y�M�3��h�����]�< ��׈��	����� �I 3�ފk��\��� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E���E�M谌���} v�MQ�M��������C����ӋU�E��M�J�E]����������������������������U��Q�M��E��HQ觫�����U��BP蘫�����M��QR艫�����E��HQ�z�������]��������������������������U��Q�M��E��HQ�G������U��BP�8������M��QR�)�������]�������������������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��E���M��B�Ћ�]���������U��Q�M��E���M��B�Ћ�]���������U��Q�M���]� ���U����M�j_h���EP�MQ�#�����j`h���UR�EP�������M���Q�UR�EP�MQ�UR�?������E��}� }	�E�������}� u	�E�    ��E�   �E��E�E��]� �����������������������������������U����M��E�    �E��HQ�M�>����U����U��E��]� ���������������U��Q�M��E��@��]����������������U��Q�M��E��@��]����������������U��Q�M��E��@��]����������������U����M��E�    �EP�M�$����M����M��E��]� ������������������U��j�hd�    P��D���3ŉE�P�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M��q����E�    �EP�MQ�������Ѕ�t�E$����U$�
�M�觞����u�E$����U$�
�P�M�蠔���E��E�    �E�Pj �M�Q�U�R诸�����]��E�;E�t�}� t�M$����E$���M(�E���U�E��M�J�E������M��N����E�M�d�    Y�M�3�������]�$ �����������������������������������������������������������������������������������U��j�hHd�    P��<���3ŉE�VP�E�d�    �M��E�P�M Q�UR�EP�MQ�U�R�M�� ����E�    �M��Z����E��EP�MQ�o������Ѕ�t�E$����U$�
�}� u�E$����U$�
�   �E�    �E�P�M(����j �M��̒�����-u)�UĉU��E�P�M(貒���   k�
�L��Uă��U��	�Eă��EċM�;M�s#�U�R�M��|����0�E�P�M(�m����L5���̋U�E��M�J�E������M�衘���E�M�d�    Y^�M�3��T�����]�$ �����������������������������������������������������������������������������������������������������U��j�h�d�    P��p���3�P�E�d�    �M��E�P�M�~����E܋M܉M��E�    �U�R��������E��E������M��@����E�    �E(�E�M��A�M�}�8�K  �U������$����M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��I�����P�M�U�  �E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�荰����@�U�E��  h`��M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�葃����P�M�U�  �E�P�M�Qjcj �UR�EP�M�Q��������U �M ��U ���ukM�d��l  �U$�J�Q  �E�P�M$��Qjj�UR�EP�M�Q�������U �M ��  h|��U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��ق����P�M�U��  �E�P�M$��Qjj �UR�EP�M�Q�2������U �M ��  �U�R�E$��Pjj �MQ�UR�E�P� ������M �U ��~  �E�P�M$��Qhn  j�UR�EP�M�Q��������U �M ��I  �U�R�E�Pjj�MQ�UR�E�P�������M �U ��E ���u�U���E$�P�  �M�Q�U$��Rj;j �EP�MQ�U�R�T������M �U ���  h���E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�茁����@�U�E�  h��j �MQ�UR�*������E�}� }�E ����U �
�kE��M$A�U$�B�Q  h���E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M�������@�U�E�  h���M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��΀����P�M�U��  �E�P�M$Qj;j �UR�EP�M�Q�*������U �M ��  h���U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��b�����P�M�U�k  �E�P�M$��Qj5j �UR�EP�M�Q�������U �M ��9  �U�R�E$��Pjj �MQ�UR�E�P�������M �U ��  �E�P�M$��Qj5j �UR�EP�M�Q�W������U �M ���   hБ�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M������P�M�U�   �E�P�M�Qjcj �UR�EP�M�Q��������U �M ��U ���u �}�E}�M��d�M���U�U��E$�M��H�B�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��������P�M�U��E ����U �
�EP�MQ�3������Ѕ�t�E ����U �
�E�M��U�P�E�M�d�    Y��]�( �I �<���,�i���G�7�t�����D�	�t���͝�y������v���>� 	
	 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��D���3�P�E�d�    �M�h  h��EP�MQ�UR�EP������h  h��M$Q�J������U�R�M�֤���E��E��E��E�    �M�Q�S������E��E������M��}���M��ҩ���E�}� u�E�   �UR�EP�������ȅ�t�  �M�y�����Rj�M�褮������u?�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M��������P�M�U�E�   �   �}�u>�E�P�M$��Qjj�UR�EP�M�Q苿�����U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P�G������M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��X�����@�U�E�MQ�UR����������t'�M�Z�����QjH�M�腭���Ѕ�t
�M������EP�MQ诜�����Ѕ�t<j �M������P�M�������E��M��:t�U��,t	�E��/u�M�k����MQ�UR�\���������t'�M�ɕ����QjH�M�������Ѕ�t
�M�/����EP�MQ��������Ѕ�t��   �M膕����Pj�M�豬���ȅ�uW�}�u�U ����M ��@�U$R�E P�MQ�UR�EP�MQ�UR�E�P�M��������P�M�U�}�u�E�   �w�}�t�}�u>�E�P�M$��Qjj�UR�EP�M�Q�z������U �M ��U$�B���M$�A�-�U�R�E$��Pjj�MQ�UR�E�P�<������M �U ��EP�MQ�������Ѕ�t'�M脔����PjH�M�诫���ȅ�t
�M�����UR�EP�ٚ�����ȅ�t<j �M�D�����R�M������E��E��:t�M��,t	�U��/u�M蕄���EP�MQ膚�����Ѕ�t'�M������PjH�M������ȅ�t
�M�Y����UR�EP�#������ȅ�t�U ����M ��  �M裓����Rj�M��Ϊ������uM�}�t�M ����E ��3�M$Q�U R�EP�MQ�UR�EP�MQ�U�R�M�������P�M�U�   �}�u>�E�P�M$��Qjj�UR�EP�M�Q觻�����U �M ��U$�B���M$�A�h�}�u/�U�R�E$��Pjj�MQ�UR�E�P�c������M �U ��3�E$P�M Q�UR�EP�MQ�UR�EP�M�Q�M��t�����@�U�E�MQ�UR����������t�M ����E ��M�U��E�A�E�M�d�    Y��]�  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M�h}  h��EP�MQ�UR�EP�V�����h~  h��M$Q��������U��BPj �MQ�UR�=������E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U��j�h�d�    P�����3�P�E�d�    �M�h�   h��EP�MQ�UR�EP�w�����h�   h��M$Q�
������U�R�M薜���E�E�E��E�    �M�Q�������E��E������M��Xu���U�R�E$��Pjj �MQ�UR�E�P�������M �U ��E �8 uj �M�6�����Q�M��ݐ���Ѓ�:t�E ����U �
�2�E�P�M$��Qj;j �UR�M�{��P�E�P�z������M �U ��E �8 uj �M�ώ����Q�M��v����Ѓ�:t�E ����U �
�/�E�P�M$Qj;j �UR�M���P�E�P�������M �U ��E�M��U�P�E�M�d�    Y��]�  ����������������������������������������������������������������������������������������������������������������������������U����M�hn  h��EP�MQ�UR�EP�f�����ho  h��M$Q��������U��BPj �MQ�UR�M������E��}� }�E ����U �
��E����M$�A�U�E��M�J�E��]�  ��������������������������������������������U��j�hd�    P�����3�P�E�d�    �M�h�  h��EP�MQ�UR�EP臿����h�  h��M$Q�������U�R�M覙���E�E�E��E�    �M�Q�#������E��E������M��hr���E�    �U�R�E�Ph�  j �MQ�UR�E�P�������M �U ��E ���u6�}�l  |�U���l  �U���}��   ~�E ����U �
�E$�M��H�U�E��M�J�E�M�d�    Y��]�  ��������������������������������������������������������������������������������U����M��E�    �E��HQ�M�����U����U��E��]� ���������������U��Q�M�j{h���EP�MQ�������U+UR�EP�V�������]� �������������������������U��Q�M��E��H$�U�
�E��]� ���������������������U����M��E�    �E��HQ�M�N����U����U��E��]� ���������������U��Q�M������]� ����������������U��Q�M��E��H �U�
�E��]� ���������������������U����M��E�    �E��HQ�M辵���U����U��E��]� ���������������U��j�hPd�    P��X���3ŉE�P�E�d�    �M��E�P�M�˖���E��M��M��E�    �U�R�H������E��E������M��o���E�P�   k���t�R�   k� ��t�Q�M�蕍���E� �E�    �M 赾���Ѕ�u+j �M ��{��� �   k�
�L�;�u�E��U����U��M �j����E��E��E��	�M����M��U�;U�s%�E�P�M �s{�����R�E�P�:�������
s�ʋM�+M�Q�U�R�M �G{��P�M������E�   �M���������t�   k� �D�Pj�M������   k� �D�P���̉e��U�R蚆���E��E�P�MQ�UR�EP�MQ�UR�EP�M������E������M�����E�M�d�    Y�M�3��b�����]� �����������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��p���3ŉE�P�E�d�    �M��E� ���] ����Au�E��E ���] �E�    �	�E���
�E��E �(�����u�}��  s�E �5��] �Ѓ��E �$hH�j(�M�Q觪�����E��}� }�U�E��M�J�E��   �U�R�M�ۓ���E��E��E��E�    �M�Q�X������E��E������M��l��j0�M������E�j �U�R�M�菂���E�   j �M��w��P�E��L�Q�   k� �L�Q�M�腊���U�R�E�P�M�躅���M�Q���̉e��U�R�Z����E��E�P�MQ�UR�EP�MQ�UR�EP�M��Κ���E������M��n}���E�M�d�    Y�M�3��"�����]�  �������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��P���3ŉE�P�E�d�    �M�h  h��EP�$�����h	  h��MQ�؛��������U蠈��E�M��I����E�    �M$��u�   ��E �D���   ��U$�T�   k��U �T��E�   ��E����E�j �M�Q�M������M����\���P�UR�E�P�M�����P�M�Q�M��{����E��U��U��E��M��g���P�S������E��}� v	�E�   ��E�    �E��E��E� �M��~����M˅�t��i����UR�EP�M�Q�M��$u��Pj�M��u��P�UR蘌�����E������M��V{���E�M�d�    Y�M�3��
�����]�  �����������������������������������������������������������������������������������������������������������U��Q�M��E��@��]����������������U��j�hHd�    P��\���3ŉE�VP�E�d�    �M��E�    jhh���EP�MQ�Ɋ�����M��7����E�    �U+U�Ũ}� ��   �E�P�M�������M���Q�UR�EP�M�Q�M�謜���E��U��U��E��M�蘯�����M���}���V�E�P�M��~����E��M��M��E��M��j���P衸�����E̍M��}��9E�w	�E�   ��E�    �UȈU��E��M��z����E� �M��n����EӅ�t��6����M�Q�M�� ����U�R�M� y���Eă��E��E������M��Qy���E�M�d�    Y^�M�3�������]� �����������������������������������������������������������������������������������������������������U��Q�M��E�P�M������M�AP�M������E��]� ���������������������U��Q�M��E���M��B$�Ћ�]���������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P�ҋE��]�  �������������������U��Q�M��E$P�M Q�UR�EP�MQ�UR�EP�MQ�U���M��P �ҋE��]�  �������������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U��Q�M��EP�MQ�U���M��P(�ҋ�]� ������������U��Q�M��EP�M���M��B,�ЋE��]� ���������������U����M��E�    �EP�M���M��B �ЋM����M��E��]� �������������U��Q�M��EP�M���M��B(�ЋE��]� ���������������U����M��E�    �EP�M���M��B�ЋM����M��E��]� �������������U����M��E��H;Mr�M��y��;Es�M��Ǚ���U��B+E;Es�M��Q+U�U�M�y��+E�E��E�;Es�M��M���+U�E��H+M;�w�M�蠍���U��B+E+E�E��M��QU+U�U�E��H;M�sj �U�R�M��n���E�;EtS�M�Q�M�賉��EEP�M�褉��EEP�q�����UR�M�Z���EP�M��}���EP�W������  �E;EwS�MQ�M��X���EP�M��L���EP�Gq�����U�R�M��4���EEP�M��%���EEP�q�����9  �E;EwS�M�Q�M������EEP�M�����EEP��p�����UR�M��ӈ��EP�M��ǈ��EP��p������   �EE;EwX�M�Q�M�蟈��EEP�M�萈��EEP�p�����UR�M��u����MM+M�P�M��a���EP�\p�����{�UR�M��G���EP�M��;���EP�6p�����E�P�M��#���EEP�M�����EEP�p�����M+MQ�M������EEP�M�����EEP��o�����U�R�M��p���E���]� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����M��} th�  hXo�EP�t�����MQ�M��r_���Ѕ�t+�EP�M��Ć���M+�Q�U�R�EP�MQ�M��{y���  �U��B;Es�M��
����M��Q+U;Us�E��H+M�M���+U�E��H+M;�w�M�������U��B+E+E�E��M;Ms*�U�R�M��:���EEP�M��+���EEP�#n�����} w�} v~�E��HM+M�M�j �U�R�M���j������tZ�M;Ms*�U�R�M��؅��EEP�M��Ʌ��EEP��m�����EP�MQ�M�誅��EP脓�����U�R�M��En���E���]� �������������������������������������������������������������������������������������������������U��j�h�d�    P��   ���3�P�E�d�    �M��E�   �E,P�M 谯���ȅ���   ���̉e��UR�����EȋEȉE��E����̉e��UR�����E��E�苝�����EЋE�P��p���Q�M��Ғ���E��U��U��E����̉e��E�P誒���E؋M؉M��E����̉e��UR茒���E��E��*������E�E�P�M��i����E���p����}����   �M Q�M,����P�M �P���P���̉�|����UR�0����E�E�E��E����̉e��UR�����E��E�谜�����E�E�P��d���Q�M�������E܋U܉U��E����̉e��E�P�ϑ���E̋M̉M��E�	���̉e��UR豑���E��E��O������EċE�P�M������E���d�����|���M��M��E��M��f���E��M��f���E� �M �|���E������M,�|���E��M�d�    Y��]�0 ��������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M�j �EP�M���l����]� ���������������������U��Q�M��E��M;Hw�UR�M���j����EP�M��U+QR�M��u����]� �������������������U��Q�M��E���M��B�Ћ�]���������U��j �EP�MQ�UR�D�����]����������������������U���   ���3ŉE��E��\����MQ�UR�_������E��E�����X����} t	�M�    �U�����U��}��  j��l���P�MQ�UR��\���P�=�������h���Q�p��$j�M�Q��[������h��� uQ���$j�U�R�[�����   ǅx���   �   �� ��l���Qj�U�R�c[������x���;�h���}Y�M�Qj�U�Rj�E�P�%_������x�������x�����x������l���Pj�M�Q�[����j�U�Rj�E�P�+[����뙋MQ�   k� �M�l���Q�U�R�(�����ٝ|����d  �}��*  j��l���P�MQ�UR��\���P蓧������`���Q�l��$j�M�Q�Z������`��� uQ���$j�U�R�Z�����   ǅt���   �   �� ��l���Qj�U�R�<Z������t���;�`���}Y�M�Qj�U�Rj�E�P��]������t�������t�����t������l���Pj�M�Q��Y����j�U�Rj�E�P�Z����뙋MQ�UR�E�P������ٝ|����   k� ��l���P��|���Q�������0�}�u��ٝ|�����}�u��ٝ|������ٝ|�����X��� t-��|���R�ck������d�����d������ �  ��d���f�
م|����M�3���z����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR��|����]����������������������U���(  ���3ŉE��E�������MQ�UR�/��������������������������} t	�M�    ����������������������  j�E�P�MQ�UR������P������������������$j�M�Q������������ u�����$j�U�R��������   ǅ����   �   �� �L�Qj�U�R�g�����������;�����}Y��0���Qj�U�Rj�E�P�p��������������������������D��Pj�M�Q������j�U�Rj�E�P訡����뙋MQ�   k� �ML�Q�U�R聡����ݝ�����t  �������1  j�E�P�MQ�UR������P�Y��������������x��$j��`���Q������������� u�����$j�U�R�׃�����   ǅ����   �   �� �L�Qj�U�R�?�����������;�����}b�� ���Qj��`���Rj�E�P�E��������������������������D��Pj��x���Q������j��x���Rj�E�P�w�����됋MQ�UR�E�P�\�����ݝ�����   k� �D�P������Q蔠�����6������u�h�ݝ�����������u�x�ݝ�������ݝ���������� t-������R�v������������������� �  ������f�
݅�����M�3��v����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR� �����]����������������������U���(  ���3ŉE��E�������MQ�UR�߃�������������������������} t	�M�    ����������������������  j�E�P�MQ�UR������P豁����������������$j�M�Q辆���������� u�����$j�U�R蟆�����   ǅ����   �   �� �L�Qj�U�R������������;�����}Y��0���Qj�U�Rj�E�P�8��������������������������D��Pj�M�Q�ʅ����j�U�Rj�E�P�y�����뙋MQ�   k� �ML�Q�U�R�φ����ݝ�����t  �������1  j�E�P�MQ�UR������P�	��������������x��$j��`���Q薅���������� u�����$j�U�R�w������   ǅ����   �   �� �L�Qj�U�R������������;�����}b�� ���Qj��`���Rj�E�P���������������������������D��Pj��x���Q蜄����j��x���Rj�E�P�H�����됋MQ�UR�E�P誅����ݝ�����   k� �D�P������Q�D������6������u��ݝ�����������u���ݝ�������ݝ���������� t-������R��g������������������� �  ������f�
݅�����M�3��[r����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} u�E�E�M�M��	�U����U��E��Q耋������t��U����-t�M����+t	�E�+   ��E���M��U����U��E��E��MQ�UR�EP�M�Q�_�����E�U�E�;u�M�U��E�M;u�}� u$�U���+u	�}����w�E���-uC�}�   �v:�,���� "   �} t	�M�   �U���-u	�E�   ���E�����E����E���-u
3�+M�M���U�U�E��]���������������������������������������������������������������������������������������U��j �EP�MQ�UR�M~����]����������������������U���$�} t	�E�     �M�M��	�U����U��E��Q�͉������t��U����-t�M����+t	�E�+   ��E���M��U����U��E��E��} |�}t�}$~�} t�M�U�3���  �   �} ~D�}u<�E����0u1�   �� �E����xt�   �� �E����Xu	�U����U��U�E����0t	�E
   �A�   �� �E����xt�   �� �E����Xu�E   �U����U���E   �E��E��	�M����M��U����0u���E�    �M��M��E�    �	�U����U��EP�M��R�֋����P�   k� ����Q�t�����E�}� t#�U�U�E�-���E��M��M�U�ʉM�렋E�;E�u�} t�M�U�3��   �E�+E܋M����+E�y�L�}� !�E��M�+�9M�r�U��E�+�3��u;E�t%����� "   �} t	�E�    �E������E�+�M���-u3�+U�U�} t�E�M���E��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�{����]����������������������U���(�} u�E��E�M�M��	�U����U��E��Q耆������t��U����-t�M����+t	�E�+   ��E���M�U����U��E�E��MQ�UR�EP�M�Q�������E�U�U�E�;u�M�U��E�M;u�U�U�u4�E���+u�}����w"r�}��w�M���-u\�}�   �rSw�}� vK����� "   �} t	�U�   �E���-u�E�    �E�   ���E������E�����E��U��2�0�M���-u3�+U�    E�U؉E���M�M؋U�U܋E؋U܋�]���������������������������������������������������������������������������������������������U��j �EP�MQ�UR�͕����]����������������������U���<V�} t	�E�     �M�M��	�U����U��E��Q茄������t��U����-t�M����+t	�E�+   ��E���M�U����U��E�E��} |�}t�}$~�} t�M�U�3�3��]  �   �} ~D�}u<�E����0u1�   �� �E����xt�   �� �E����Xu	�U����U��U�E����0t	�E
   �A�   �� �E����xt�   �� �E����Xu�E   �U����U���E   �E��E��	�M����M��U����0u���E�    �E�    �M��M��E�    �E�    �E� �	�U����U��EP�M��R聆����P�   k� ���Q�Xo�����E��}� t@�U܉UԋE��E؋M�����M��E�RP�U�R�E�P�֖���ȋ��E����M܉u�냋U�;U�u�} t�E�M�3�3���   �U�+U�E���+щU�y�   �}� Y�E���M�+ȋE�M̉EЋM�;M�r<w�U�;U�r2�E���M�+ȋu��E�RPVQ�,a���EĉUȋU�;U�u�E�;E�t,�o���� "   �} t	�M�   �E������E������E�+�U���-u3�+Eܹ    M��E܉M��} t�U�E���E܋U�^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����l���E��uH���   �� ��U��}� t�E�P�v�����E��E��U���]�����������������U���$�E�    �E+E�E�M+M�M��} u�H���   �� ��E��l���E���M�Q�U��E��M܃}� ui�U�;U�}�E�E���M��M�U�R�EP�MQ�PP�����E�}� u(�U�;U�t �E�;E�}	�E�������E�   �M�M���U�U��E��E��M�M�Q�U�R�EP�M�Q�URh   �E�Pj ��n���� �E��}� u�
����    �E�����	�M����M��E���]���������������������������������������������������������������������������U���3�f�E�3�f�M�j�U�Rj"�F���   k��P�-D�����   k� �D���0u	�E�   �I�   k� �D���1u	�E�   �(�   k� �D���2u	�E�   ��E�    �M��M�U�U��E���]���������������������������������������������������U���l���3ŉE�VW�} t�} u3��@  �E���u�} t3ҋEf�3��!  �} u�M�Q�#������   ���}��UЉU�E�x t�} t�Mf��Ef��   ��  �M�yt,�U�zt#hP�h�Yj j^h��j��D������u̋M�9 ��   �   �� �E�M�	��U�zv6�} t	�E�   ��E�    �E�P�MQj�URj	�E�Q� ��u�U�    袊��� *   ����(  �E�     �M�A�  �U��E��M����U�D
�Mσ��   ��#���   �E�M;Hs�   k� �M�U��������   �h�E�xv;�} t	�E�   ��E�    �M�Q�UR�E�HQ�URj	�E�Q� ��u$�U�B��u�M�    �̉��� *   ����U�U�B�M�K�} t	�E�   ��E�    �E�P�MQj�URj	�E�Q� ��u�|���� *   �����   _^�M�3���a����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��� �E+E���E�M+M���M��E�    �} u�B���   �� ��E��	�M�Q�U��}� ui�E�;E�}�M�M���U��U�E�P�MQ�UR��   ���E�}� u(�E�;E�t �M�;M�}	�E�������E�   �U�U���E�E��M��M��G�U�R�EP�M�Q�URh   �E�P�sj�����E��}� u�̇���    �E�����	�M����M��E���]�����������������������������������������������������������������������������U��Q��E���E�M���M�U���U�} ~7�E��U�;�t%�M��E�;�}	�E�������E�   �E���3���]�����������������������������U����E+E���E�M+M���M��E������E�    �} u��@���   �� ��E��	�M�Q�U�}� u)�E�;E�w�M���Q�UR�EP�dI�����M�M��   jgh$�j�U�R�<�����E��}� ��   �E�P�M�Q�U�R�EPh   �M�Q��y�����E��}� u/j j �U�R�EPh   �M�Q��y�����E��}� u�E�����0�E�    �	�U����U��E�;E�s�M�M�f��E��Mf�A�ك}� tj�U�R��M�����E���]����������������������������������������������������������������������������������������������U����E�Pj�MQj� ��u	�E�    ��U��U�f�E���]�����������������������������U��EP�M+M��Q�URj� �E]����������������U��Qf�Ef�E��M����  u�_�U�z u*�E=   }�M��A|�U��Z�E�� f�E��,j�M�Qj�URh   �E�HQ�'x������uf�Uf�U�f�E���]������������������������������������������������U��Qf�Ef�E��M����  u�_�U�z u*�E=   }�M��a|�U��z�E�� f�E��,j�M�Qj�URh   �E�HQ�ww������uf�Uf�U�f�E���]������������������������������������������������U����E+E�E�M+M�M��E������} u�n=���   �� ��E��na���E���M�Q�U�E��M��}� u*�}� u$�U�;U�w�E�P�MQ�UR��E�����E��E��ej�M�Qj j �U�R�EPh   �M�Qj �[u����$�E��}� t7�U��U�E�;E�)j�M�Q�U�R�EP�M�Q�URh   �E�Pj �u����$�E��]������������������������������������������������������������������U����E��M��E�    �	�U����U��E��Q�t������t��U����-u�E�   �M����M���U����+u	�M����M��U����nt�M����N��   �E����E��M����at�E����Au�U����U��E����nt�U����Nt�M��U��E�    �d�E����E��M��M��E�   �U����(uC�M����M��U��P���������u�M����_u�׋E����)u�U����U��E��E��} t�M�U����  �E����it�U����I�"  �M����M��U����nt�M����Nu�E����E��M����ft�E����Ft�U��E��E�    �   �M����M��U��U��E���E�M����it�E����I��   �U����U��E����nt�U����Nul�M����M��U����it�M����IuM�E����E��M����tt�E����Tu.�U����U��E����yt�U����Yu�M����M��U��U��} t�E�M���   �U����0uw�   �� �U��
��xt�   �� �U��
��XuO�M����M�U����.u	�M���M�U��P��z������u�M���M���U����U��E���E��	�M���M�U�E���E��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���l���3ŉE�V�E�    kE	�E�}-~�E-   �   k� �E�    �   �� �U�
    �E�    ��E���E�E�   �M���0u���E�    ��E���E�E�   �M�R�r�������tD�E�;E�M���0�EȈT̋Mȃ��M���   k� �M����   k� �E�뙋M�1��J���   k� ��
;�u	�M���M�}� u>��U���U�E�   �E���0u!�   k� �M����   k� �E�����M���M�E�   �U�P蟃������tB�M�;M8�U���0�MȈD̋Uȃ��Uȸ   k� �U�
���   k� �M�뛋U;U�}I�E�E��M��T̃�|�E��Lˀ��U��LˋE�Eȹ   k� �E����   k� �U��	�Eȃ��Eȃ}� ~-�M��T˅�u!�   k� �U�
���   k� �M��ă}� u$�UȉU��Eȃ��Eȃ}�.s��Yt���M��D� �}� ��  �E�    �Eș�	   ���	   +E��E���	   ����u	�E�    ��E�   �U��U���E����E��M����M��U�;U�}J�E���	   ����u�Uă��UċE��L̋UċE����MċUk�
�M��T�MċU��뜋E���et�U���E��   �M�M��U���U�E���+t�U���-t	�E�+   ��M��U��E���E�M��M��E�    �E�    ��U���U�E�   �E�Q�`�������t�}� ��}kU�
�E��T
ЉU����E���-u�M��ىM��   k� �M�U��   k� �E��}� u�M��M�}� u�E�    �} t�}� t�U�U���E�E��M�U���E�^�M�3��pR����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���d���3ŉE�V�E�    kE�E�}#~�E#   �   k� �E�    �   �� �U�
    �E�    ��E���E�E�   �M���0u���E�    ��E���E�E�   j�M�R�   k� ��X�Q�3W�����E��}� tL�U�;U �E�-X��MԊ�p��T؋Eԃ��E���   k� �E����   k� �U��{����E�0�sE���   k� � �;�u	�U���U�}� u>��E���E�E�   �M���0u!�   k� �U�
���   k� �M�����U���U�E�   j�E�Q�   k� X�P�CV�����E��}� tH�M�;M>�U���X��EԊ�p��L؋Uԃ��UԸ   k� �U�
���   k� �M�뀋U;U�}I�E�E��M��T؃�|�E��L׀��U��L׋E�EԹ   k� �E����   k� �U��	�Eԃ��Eԃ}� ~-�M��Tׅ�u!�   k� �U�
���   k� �M��ă}� u$�UԉU��Eԃ��Eԃ}�$s���n���M��D� �   k� �M����   k� �E��}� ��  �E�    �Eԙ�   ���   +E��E���   ����u	�E�    ��E�   �U��U���E����E��M����M��U�;U�}L�E���   ����u�UЃ��UЋE��L؋UЋE����MЋU�����M��T�MЋU��뚋E���pt�U���P��   �M�M��U���U�E���+t�U���-t	�E�+   ��M��U��E���E�M��M��E�    �E�    ��U���U�E�   �E�Q�{������t�}� ��}kU�
�E��T
ЉU����E˃�-u�M��ىMĺ   k� �M�Uĸ   k� �E��}� u�M��M�}� u�E�    �} t�}� t�U�U���E�E��M�U���E�^�M�3��L����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�E��   �� �U��
%�  =�  u?�   �� �U��
��u�   k� �E����u	�E�   ��E�   f�E��]�[�   �� �E�������u�   k� �M����t/�   �� �M����  u	�E�������E�����f�E���3���]������������������������������������������������������������U��   k� E]�����������������U��   �� E]�����������������U���(V�E�E�   �� �U��
%�  ��f�E��M����   uB�   �� �E����u�   k� �M����u	�E�   ��E�   f�E��i  �'�E���u�M�Q�nk����f�E��U���~3��@  �} ~T�E���   +�;MD�   �� �E���� �  t�����]��	���]��U�E���   ��  ��  �E���;E}<�   �� �U��
%����M�M����   �� �M�f�����  �  �   �� �E���� �  f�M�   �� �E�����ɀ   �   �� �E�f��M��U�D
��E�}�|�} |0�   �� �U�f�E�f�
�   k� 3��M�f�3��  �  f�Uf�U�3�f�E��M����h�U��t	�E�   ��E�    �   k� �U��
E�f�E��   �� �   k� �U�u�f�f��   �� 3��M�f��U���f�U��E���f�E��M�����   �U��t	�E�   ��E�    �   k� �U��
�M��   +ы���E�f�E��   k� �U��
�M����   �� �U��
�M��   +����º   k� �U�f�
�   �� �M�f�f�M�f��   �� �M�f��   �� �E��M��и   �� �M�f��U�� �  �E�= �  un�   k� �E����tZ�   k� �M�f�f��f�U�   k� �U�f�E�f�
�M����  u$�   �� �E�f�f���   �� �E�f��.�   �� �U��
�M�;�u�   k� �M����u3�����^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���<V�E�]܃} u�  �E�P�M�Q�T����f�E��U�����   �E���t �   k� UR�X����f�E��E����   k� �E�E��u�M���t6�UR� 5�����0�� �  �   k� MQ�5������� �  ;�u�4j�i3�����   k� �U���
�}~�   �� �M�����  �U�����  �E�   �E�    �E�;E��  �M��U���]��E�   �E�P�M�Q�S����f�E��U���~
�|  �r  �E���u-�M��U�E���E���;E}�M��U���\��G  �=  �E��M�+��EԋU���9U���   �E��������D��   �E��E�M���M�U�;U}�E�M����������D{�ًU��9U�}�E���E���M�;Mu	�U���U��	�E���E�M�;M�}�U�E�M�u�D�����ڋU��E�E�����]�~  �M�;M�#�E��������D{�U��U��E����E��S  �M��U���E�]ЋE��M�E����E���������Dzf�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E��M����������Dz��  �U��E���]�MQ�U�R�Q�����E�+E��M�;���   �U�E�+E�+�R�MQ��1�����U�R�EP�R�����M��U���e�]̋E��M�E����E���������DzM�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E����E�u	�E�   �$�M��U�D���]܍E�P�M�Q��P�����U��U��   �E���;Eu
�   �   �M��U���]�E��M��R�E�P�P����j�M��U��P��0�����M�Q�U��E��Q�Q�����E�U��E�$��]�M��M��E��������D{�E�]���U��E���]��E��]܍M�Q�U�R�P�����E����E��D����E^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}3�U��E����������D{�M��UQ���$�EP�MQ�&����뼋E��]�������������������������U����} u���b  �]  �}t2�   k� �U�
��������D{�   �� �M���������Dz�   k� �M��  �  �}t�   ��E���������Dz,�   k� �   �� �M��U��]��E���   ��   �   k� �   �� �E��M��]��   ��E��]��   k��E���������D{�M�Q��-�����E��U�����M�f��   k� �E�M�$�   �� �E�������Dz�E��E��]��E��'�%�   k� �   �� �M��E��E��]��E��]��������������������������������������������������������������������������������������������������������U����} u�  �   k� MQ��O����f�E��U���|<�E���u�   k� �E�����M���u�   k� �M����.  �U�U��E�M���U�E�M���U�   k� �U�
�]��EP�MQ�U�R����������$�EP�M�Q�������}~�   �� �E��E��]��E������]��E�Q�$�MQ�UR�l�����E�   ��E����E�M�;M}~�UR�EP�M�Q�K�����U�R�EP�M�Q�UR�E�P���������$�MQ�U�R�������E�P�MQ�UR�EP�M�Q������UR�E�P�MQ�UR�������r����E��]���������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}<�UR�E��M�����$�V�����U��E���M��U����������Dz�볋E��]��������������������������������U��E��P�MQ�UR��$�����E]������������������U���0���3ŉE��} ��   �   k� �U�
�M�   k� �\�   k� �L�Q�M����f�E��U���|S�E���u
j�(�����   k� �   k� �E�D���M���~�}~�   �� �E����E�  �   k� �E����E�   �E�    ��M���M�U���U�E�;E�L  �	�M���M�}�}\�U�U�;U}=�E�E�M����������D{&�U�U�E���M�M��\��U�U�E������M����\���E�   �땺   k� �D���������Dz
��   �   �E�    �   k� �D��]؍E�P�M�Q�H����j�U�R�l(�����E�P�M�Q�?I�����E��$�UR�EP������   k� �D��e��]��E�Q�$�EP�MQ�j�����U܃��U܋E�;E�}$�M܋U��D���\��E��D����������Dz��������E�M�3��8����]�����������������������������������������������������������������������������������������������������������������������������������������������������������U����} t�} u�  �   k� �U�
��������D{�   �� �M���������Dz'�   k� �MQ��$�UR�EP�������   �M�M�U�E���M��UR�EP�M�Q�F�����   k� �MQ��$�UR�EP�[�����E�   �	�M����M��U�;U}_�E��M����������D{K�U�R�EP�M�Q�������U��EQ���$�MQ�U�R�������EP�M�Q�UR�EP�����됋E��]�����������������������������������������������������������������������������������������U����E��'  ���E��E��]��E�Q�$�UR�EP���������$�MQ�UR�9�����E��'  ���U��E��]��E�Q�$�UR�EP������E��]�������������������������������������U����E�]�} �m  �}t�E�P�M�Q�~D����f�E��U���u�   k� �U�E��
�5  �E���~&�   k� �E�E���   �� �U���
�  j�E�P�|$�����M�Q�U�R�OE�����   k� �U�E��
�E�e��   �� �M�3���   �   �� �M��]�   �� UR�E�P�C����j�   �� MQ��#�����U�R�   �� EP��D�����   �� �E�U�$
�   ���M��}~(�   ��E���������D{�   k��E�����}~�   ��U���
�E��]������������������������������������������������������������������������������������������������������U����} u��  �   k� MQ�=F�����Ѕ�}�   k� �U�
�x^����z>�   k� �U�
�x^����zj�!�����   k� �U���
�P  �E�E��M�U���E��M�U����E��   k� �E��]��}~�   �� �E��U�
�]��E����$�X	 �������]��E�Q�$�EP�M�Q������E�   ��U���U�E�;E��   �M�Q�UR�E�P���������$�MQ�U�R������E�P�MQ�UR�EP�M�Q������U�R�EP�M�Q�UR�E�P����������$�MQ�U�R�������E�P�MQ�U�R�EP�M�Q������M����U�R�EP�M�Q�UR�EP������E��]�������������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}5�U��E����������D{!�M��U����Q�$�EP�MQ�����뺋E��]�����������������������U���8���3ŉE��} t�   k� �U�
��������Dzj�EP�������   �} ~Q����$j�M�Q�������U�ډUh��j�E�P�o�����M��t�U�Rj�E�Pj�MQ������U���Uu�,�E�Pj�M�Q�1�����U�Rj�E�Pj�M�Q�������j�UR�������]��E���������D{&�E���������D{�����E�������Dz��V��� "   �} t�E����U�
�EȋM�3��D/����]����������������������������������������������������������������������������������������U����E�E��   k��E�����  ���  ug�   k��M����uA�   ���M����u/�   �� �M����u�   k� �U��
��u	�E�   ��E�   f�E��   ��   k��E�������u8�   ��E����u&�   �� �E����u�   k� �M����t.�   k��U��
%�  u	�E�������E�����f�E���3���]������������������������������������������������������������������������������U��   k� E]�����������������U��   k�E]�����������������U���0V�E�E�   k��E�����  ��f�M��U����  ug�   k��U��
��uA�   ��U��
��u/�   �� �U��
��u�   k� �E����u	�E�   ��E�   f�E���  �'�U���u�E�P�/0����f�E��M���~3���  �} ~T�U���  +�;ED�   k��E���� �  t�h����]��	�h��]ЋU�E���   �m  �h  �E���;E}=�   k��E��������U�U��ʸ   k��E�f�����%  �   �   k��E���� �  f�M�   k��M�������   k��E�f��M��U�D
��E�}�|�} |Q�   k��E�f�M�f��   ��3��M�f��   �� 3��M�f��   k� 3ɋU�f�3��}  �x  f�Ef�E�3�f�M���U���f�U��E������   �M��t	�E�   ��E�    �   k� �M��U�f�U��   �� �   k� �M�u�f�f��   ��   �� �E�u�f�f��   k��   ��U�u�f�f�
�   k�3��M�f��L����U���f�U��E����)  �M��t	�E�   ��E�    �   k� �M���E��   +���U�f�U��   k� �E���M����   �� �M���M��   +����и   k� �E�f��   �� �U��
�M����   ��U��
�M��   +����º   �� �M�f��   ��E���M����   k��E���M��   +����и   ���M�f��   k��M�f�f�M�f��   k��E�f��   k��E��M��и   k��E�f��M�� �  (�U�� �  ��   �   k� �U��
����   �   k� �E�f�f��f�M�   k� �M�f�U�f��E�%��  ��   �   �� �U�f�
f��f�E�   �� �U�f�E�f�
�M����  uX�   ��E�f�f��f�M�   ��E�f�M�f��U����  u$�   k��U�f�
f���   k��M�f��S�   k��M���E�;�u<�   ��U��
��u*�   �� �U��
��u�   k� �E����u3�����^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���PV�E�]Ѓ} u�  �E�P�M�Q�@����f�E��U�����   �E���t �   k� UR�h3����f�E��E����   k� �E�E��u�M���t6�UR�%�����0�� �  �   k� MQ�f%������� �  ;�u�4j�Y�����   k� �U�x��
�}~�   �� �M�����  �U�����  �E�   �E�    �E�;E��  �M��U���]��E�   �E�P�M�Q�?����f�E��U���~
�|  �r  �E���u-�M��U�E�ʋE���;E}�M��U���\��G  �=  �E��M�+��E؋U���9U���   �E��������D��   �E��E�M���M�U�;U}�E�M����������D{�ًU��9U�}�E���E���M�;Mu	�U���U��	�E���E�M�;M�}�U�E�M�u�D�����ڋU��E�E�����]�~  �M�;M�#�E��������D{�U��U��E����E��S  �M��U���E�]ȋE��M�E����E���������Dzf�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E��M����������Dz��  �U��E���]�MQ�U�R�=�����E�+E��M�;���   �U�E�+E�+�R�MQ�"�����U�R�EP�qL�����M��U���e�]��E��M�E����E���������DzM�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E����E�u	�E�   �$�M��U�D���]ЍE�P�M�Q��<�����U��U��   �E���;Eu
�   �   �M��U���]�E��M��R�E�P�<����j�M��U��P�!�����M�Q�U��E��Q�\K�����U��E�E�$��]�M��M��E��������D{�E�]���U��E���]��E��]ЍM�Q�U�R�<�����E����E��D����E^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}5�U��E����������D{!�M��U�����$�EP�MQ�H����뺋E��]�����������������������U���V�} u���P  �K  �}t2�   k� �U�
��������D{�   �� �M���������Dz�   k� �M��   ��   �}t�   ��E���������Dz&�   k� �   �� �M�u���   �   �   k� �   �� �U�u���]�   ���M��]��   k��M���������D{�U�R�	�����E��E�����U�f�
�   k� �U�E��$
�   �� �M�������Dz
�E��E��!��   k� �   �� �U�
�E�M�^��]��������������������������������������������������������������������������������������������������������U����} u�  �   k� MQ�X+����f�E��U���|<�E���u�   k� �E�����M���u�   k� �M�h���(  �U�U��E�M���U�E�M���U�   k� �U�
�]�EP�MQ�U�R�F�����ؤ�$�EP�M�Q�9(�����}~�   �� �E�E���]����u���$�MQ�UR��(�����E�   ��E����E��M�;M}~�UR�EP�M�Q�F�����U�R�EP�M�Q�UR�E�P�t(�������$�MQ�U�R�BE�����E�P�MQ�UR�EP�M�Q�C(�����UR�E�P�MQ�UR�E�����r����E��]���������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}<�UR�E��M�����$�V������U��E�ЋM��U����������Dz�볋E��]��������������������������������U��E��P�MQ�UR�������E]������������������U���@���3ŉE��} ��   �   k� �U�
�M�   k� �\ܺ   k� �L�Q�q(����f�E��UЅ�|S�EЃ�u
j�	�����   k� �   k� �E�D���MЅ�~�}~�   �� �E����E�  �   k� �E����E�   �E�    ��Mԃ��MԋU؃��U؋E�;E�E  �	�M؃��M؃}�}\�U�U�;U}=�E�E؋M����������D{&�U�U؋E���M�M��\�܋U�U؋E������M����\���E�   �땺   k� �D���������Dz
�   �   �E�    �   k� �D��]��E�P�M�Q�14����j�U�R�*�����E�P�M�Q�C���E��$�UR�EP�B�����   k� �D��e����$�EP�MQ��A�����Ũ��ŰE�;E�}$�M̋U��D���\�ԋE��D����������Dz��������E�M�3������]��������������������������������������������������������������������������������������������������������������������������������������������������U����} t�} u�   �   k� �U�
��������D{�   �� �M���������Dz)�   k� �M����$�UR�EP�#������   �M�M�U�E�ЉM��UR�EP�M�Q�A�����   k� �M����$�UR�EP�"�����E�   �	�M����M��U�;U}a�E��M����������D{M�U�R�EP�M�Q�@�����U��E�����$�MQ�U�R�U"�����EP�M�Q�UR�EP�j@����뎋E��]�����������������������������������������������������������������������������������U����E�]��E����$�EP�MQ�"�����E��]���������������������U����E�]��} �  �}t�E�P�M�Q�1����f�E��U���u�   k� �U�E��
�a  �E���~&�   k� �E�E���   �� �U���
�3  j�E�P������M�Q�U�R�?�����   k� �U�E��
�E�e�   �� �M��   ����   �}��   �   �� �M���������D��   �   �� �E��]�   �� MQ�U�R�0����j�   �� EP������M�Q�   �� UR��>�����   �� �M�E�$�   ��E��}~(�   ��U�
��������D{�   k��U���
��}~�   ���M����E��]��������������������������������������������������������������������������������������������������������������������������U����} u�  �   k� MQ��!�����Ѕ�}�   k� �U���
����Au:�   k� �U���
����Auj�������   k� �U�x��
�L  �E�E��M�U�ʉE��M�U��ʉE��   k� �E��]�}~�   �� �U�E��
�]���E��$��  ��������$�EP�M�Q�v�����E�   ��U���U��E�;E��   �M�Q�UR�E�P�<�����Ȥ�$�MQ�U�R�7�����E�P�MQ�UR�EP�M�Q�������U�R�EP�M�Q�UR�E�P���������$�MQ�U�R�;�����E�P�MQ�U�R�EP�M�Q������M����U�R�EP�M�Q�UR�EP�b�����E��]���������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}7�U��E����������D{#�M��U�������$�EP�MQ�k:����븋E��]�������������������������������������U���l���3ŉE��} t�   k� �U�
��������Dzj�EP��������   �} ~�����$j�M�Q�5������U�ډUh�j�E�P�Z:�����M��t�U�Rj�E�Pj�MQ������U���Uu�,�E�Pj�M�Q�:�����U�Rj�E�Pj�M�Q������j�UR�5�����]��E���������D{&�E��h�������D{�h����E�������Dz� 8��� "   �} t�E����U�
�E��M�3��r����]��������������������������������������������������������������������������������������U��EP�n����]����������������U��   k� E]�����������������U��   k�E]�����������������U��EP�MQ�9����]������������U���PV�E�]Ѓ} u�  �E�P�M�Q�@����f�E��U�����   �E���t �   k� UR�*"����f�E��E����   k� �E�E��u�M���t6�UR�x�����0�� �  �   k� MQ�[������� �  ;�u�4j�������   k� �U����
�}~�   �� �M�����  �U�����  �E�   �E�    �E�;E��  �M��U���]��E�   �E�P�M�Q�u?����f�E��U���~
�|  �r  �E���u-�M��U�E�ʋE���;E}�M��U���\��G  �=  �E��M�+��E؋U���9U���   �E��������D��   �E��E�M���M�U�;U}�E�M����������D{�ًU��9U�}�E���E���M�;Mu	�U���U��	�E���E�M�;M�}�U�E�M�u�D�����ڋU��E�E�����]�~  �M�;M�#�E��������D{�U��U��E����E��S  �M��U���E�]ȋE��M�E����E���������Dzf�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E��M����������Dz��  �U��E���]�MQ�U�R�=�����E�+E��M�;���   �U�E�+E�+�R�MQ�7�����U�R�EP������M��U���e�]��E��M�E����E���������DzM�U��U�E���E�M�;M}*�U�E�M�u���\���U�E�D����������D{�ŋM�U���\���E����E�u	�E�   �$�M��U�D���]ЍE�P�M�Q�<�����U��U��   �E���;Eu
�   �   �M��U���]�E��M��R�E�P�o<����j�M��U��P�(�����M�Q�U��E��Q������U��E�E�$��]�M��M��E��������D{�E�]���U��E���]��E��]ЍM�Q�U�R��;�����E����E��D����E^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}5�U��E����������D{!�M��U�����$�EP�MQ�����뺋E��]�����������������������U���V�} u���P  �K  �}t2�   k� �U�
��������D{�   �� �M���������Dz�   k� �M��   ��   �}t�   ��E���������Dz&�   k� �   �� �M�u���   �   �   k� �   �� �U�u���]�   ���M��]��   k��M���������D{�U�R�������E��E�����U�f�
�   k� �U�E��$
�   �� �M�������Dz
�E��E��!��   k� �   �� �U�
�E�M�^��]��������������������������������������������������������������������������������������������������������U����} u�  �   k� MQ�����f�E��U���|<�E���u�   k� �E�����M���u�   k� �M����(  �U�U��E�M���U�E�M���U�   k� �U�
�]�EP�MQ�U�R������ؤ�$�EP�M�Q������}~�   �� �E�E���]����u���$�MQ�UR�)�����E�   ��E����E��M�;M}~�UR�EP�M�Q������U�R�EP�M�Q�UR�E�P���������$�MQ�U�R�l�����E�P�MQ�UR�EP�M�Q������UR�E�P�MQ�UR� �����r����E��]���������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}<�UR�E��M�����$�v�����U��E�ЋM��U����������Dz�볋E��]��������������������������������U��E��P�MQ�UR�,������E]������������������U���@���3ŉE��} ��   �   k� �U�
�M�   k� �\ܺ   k� �L�Q�3����f�E��UЅ�|S�EЃ�u
j��������   k� �   k� �E�D���MЅ�~�}~�   �� �E����E�  �   k� �E����E�   �E�    ��Mԃ��MԋU؃��U؋E�;E�E  �	�M؃��M؃}�}\�U�U�;U}=�E�E؋M����������D{&�U�U؋E���M�M��\�܋U�U؋E������M����\���E�   �땺   k� �D���������Dz
�   �   �E�    �   k� �D��]��E�P�M�Q�4����j�U�R��������E�P�M�Q�H���E��$�UR�EP�9�����   k� �D��e����$�EP�MQ������Ũ��ŰE�;E�}$�M̋U��D���\�ԋE��D����������Dz��������E�M�3��^����]��������������������������������������������������������������������������������������������������������������������������������������������������U����} t�} u�   �   k� �U�
��������D{�   �� �M���������Dz)�   k� �M����$�UR�EP�S������   �M�M�U�E�ЉM��UR�EP�M�Q������   k� �M����$�UR�EP������E�   �	�M����M��U�;U}a�E��M����������D{M�U�R�EP�M�Q������U��E�����$�MQ�U�R������EP�M�Q�UR�EP������뎋E��]�����������������������������������������������������������������������������������U����E�]��E����$�EP�MQ�������E��]���������������������U����E�]��} �  �}t�E�P�M�Q��0����f�E��U���u�   k� �U�E��
�a  �E���~&�   k� �E�E���   �� �U���
�3  j�E�P�N������M�Q�U�R�������   k� �U�E��
�E�e�   �� �M��   ����   �}��   �   �� �M���������D��   �   �� �E��]�   �� MQ�U�R��/����j�   �� EP�������M�Q�   �� UR������   �� �M�E�$�   ��E��}~(�   ��U�
��������D{�   k��U���
��}~�   ���M����E��]��������������������������������������������������������������������������������������������������������������������������U����} u�  �   k� MQ������Ѕ�}�   k� �U���
����Au:�   k� �U���
����Auj�$������   k� �U����
�L  �E�E��M�U�ʉE��M�U��ʉE��   k� �E��]�}~�   �� �U�E��
�]���E��$������������$�EP�M�Q������E�   ��U���U��E�;E��   �M�Q�UR�E�P������Ȥ�$�MQ�U�R������E�P�MQ�UR�EP�M�Q�,�����U�R�EP�M�Q�UR�E�P���������$�MQ�U�R������E�P�MQ�U�R�EP�M�Q�������M����U�R�EP�M�Q�UR�EP������E��]���������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �	�E����E��M�;M}7�U��E����������D{#�M��U�������$�EP�MQ�����븋E��]�������������������������������������U����E�$���  ��]�����������U���l���3ŉE��} t�   k� �U�
��������Dzj�EP��������   �} ~�����$j�M�Q�E������U�ډUh�j�E�P�F�����M��t�U�Rj�E�Pj�MQ�������U���Uu�,�E�Pj�M�Q������U�Rj�E�Pj�M�Q������j�UR�9�����]��E���������D{&�E���������D{�����E�������Dz�@!��� "   �} t�E����U�
�E��M�3�������]��������������������������������������������������������������������������������������U���V�   �� �M��� �  f�U��   f�E��   �� �U�
���E��   �� �Uf�E�f�
�M��u�   k� �M����e  �   �� �M���u:�   k� �   �� �E�uf�f��   k� 3ɋUf��E���f�E��f�M�f��f�M��   �� �E����   }W�   �� �E���   k� �U���Ⱥ   �� �Ef��   k� �Ef�f��   k� �Uf���f�E�f��f�E��   �� �U�
=   |W�   k� �E����   �� �E���ʸ   k� �Ef��   �� �Uf�
f��   �� �Uf�
뇸   �� �M����   �� �Mf��   �� �E��M�и   �� �Mf�f�E�^��]�����������������������������������������������������������������������������������������������������������������������������������������������U��E��t�!��� !   ��M��t���� "   ]��������������������U����E�E��   �� �U��
%�  ��f�E��M����   uB�   �� �E����u�   k� �M����u	�E�   ��E�   f�E��Z  �1�   �� �M�������u�   k� �U��
��u3��'  �M���   +��E+�f�U��M���3��  ��   �U���|B�   �� �M���� �  �   �� �M�f��   k� 3ɋU�f�����   �   �E���f�E4�f�M�f�U�f��f�U��E���T��U��J�M�#�f�M��U���T��M��U��B3��M���T��M�f�Q�U���~*�   k� �U��
�M��f�M��   k� 3ɋU�f��E���t	�E�������E�    f�E��]��������������������������������������������������������������������������������������������������������������������������������U����E�E��   �� �U��
%�  ��f�E��M����   uG3ҋEf��   �� �U��
��u�   k� �E����u	�E�   ��E�   f�E��j�h�U����E�P�:����f�E��M���>�   �� �E��������� ?  �   �� �E�f��M���~�Uf�
�����
3��Mf�3���]�����������������������������������������������������������U���V�   k��U�
% �  f�E��   f�M��   k��M����U��   k��Uf�E�f�
�M��u<�   ��E���u*�   �� �E���u�   k� �M����y  ��E���f�E��   k��E���un�   ��   k��E�uf�f��   �� �   ��U�uf�f�
�   k� �   �� �M�uf�f��   k� 3ҋEf��t����f�M�f��f�M��   k��M�����   �   k��U�
��   ��U�
����   k��Uf�
�   ���M���   �� �M���й   ��Ef��   �� �U�
��   k� �M���¹   �� �Uf�
�   k� �Uf�
f��   k� �Mf������f�U�f��f�U��   k��U�
�� ��   �   k� �E����   �� �E���ʸ   k� �Ef��   �� �U�
���   ��U�
����   �� �Mf��   ��E����   k��U���Ⱥ   ��Ef��   k��Ef�f��   k��Uf������   k��U�
���   k��Mf��   k��M��U���   k��Mf�f�E�^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�E��   k��E�����  ��f�M��U����  ug�   k��U��
��uA�   ��U��
��u/�   �� �U��
��u�   k� �E����u	�E�   ��E�   f�E��  �V�   k��M�������u?�   ���M����u-�   �� �M����u�   k� �U��
��u3��  �M��3  +��E+�f�U��M���3��  �  �U���5|b�   k��U��
% �  �   k��M�f��   ��3��M�f��   �� 3��M�f��   k� 3ɋU�f�����  �  �E���f�Ed�f�M�f�U�f��f�U��E������U��J�M�#�f�M��U������M��U��B3��M������M�f�Q�U��U��}�t`�}�t0�}�t�|�   ���M���E��f�E��   ��3ҋE�f��   �� �U��
�M��f�M��   �� 3��M�f��   k� �M���E��f�E��   k� 3��M�f��U���t	�E�������E�    f�E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�E��   k��E�����  ��f�M��U����  ul3��Mf��   k��M����uA�   ���M����u/�   �� �M����u�   k� �U��
��u	�E�   ��E�   f�E��l�j�M����U�R�{�����f�E��E���@�   k��E����������?  �   k��U�f��E�-�  �Mf������
3ҋEf�3���]�����������������������������������������������������������������������������������U���EP�MQ������]�����������U��EP�MQ�{����]������������U��SV��څ�t��t�U��tW�̋�����F�^�2_^[]� ��������������U��QS�ډM�VW��tM3�93~G3����    �K�E��9�|�����u�D9U��<����t�t9�EP�l�����F��;3|Ëu3��ƅ�t`�@G��u���tT�>����u�~����u�~����u	�~����t�EWVP��������F�|0�����t�EWVP��������vO��u�_^[��]� ���������������������������������������������������������������U��QS�ډM�V3�93~AW3��K�E��9�|�����u�D9U��<����t�t9�EP�h�����F��;3|�_^[��]�������������������������u�U��� PRSVW�Ej P�h�����_^[ZX��]�����������̀=�� uj jj j j ��������P�r�����������������������������jjj j j ���������������������U����P� ]����������������U��Q���P� �E��}� t�U�j������jj �s�����������]����������������������U��Q�E�    ���P� �E��MQ� ����E���]�����������������U��Qh�   h��jjj �������E��E�P� �h��h��d��}� u�   ��U��    3���]���������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �����E�    �EP�T   ���E��E������   �����ËE�M�d�    Y_^[��]��������������������������������������U����h�P� �E��d�Q� �E��U�;U�r�E�+E�����s3���   j�M�Q�������E�U�+U���9U���   �}�   s�E�E���E�   �M�M�M��U�;U�r"j}h��j�E�P�M�Q�h������E�}� u:�U���U��E�;E�r%h�   h��j�M�Q�U�R�2������E�}� u3��Q�E�+E����M���U��E�E��M�Q� �h��UR� �M���U����U��E�P� �d��E��]����������������������������������������������������������������������������������U��Q�EP��������u	�E�������E�    �E���]����������������������U���  ���j�s������EP�=������=�� u
j�T�����h	 ��������]���������������������������U���$  j�(�����t�   �)�������������5���=��f���f���f���f�|�f�%x�f�-t������E ����E����E������������  ���������	 ����   ���   �   k� ǂ��   �   k� ����T��   �� ����L�hХ�������]������������������������������������������������������������������������������U��j����]�����U���  j�������t�M�)�������������5���=��f���f���f���f�|�f�%x�f�-t������E ����E����E������������������	 ����   ���   �   k� �E����hХ�������]���������������������������������������������������������������U���   j������t�M�)�������������5���=��f���f���f���f�|�f�%x�f�-t������E ����E����E������������������	 ����   �} v�} u�E    �}v	�M���M�U������   k� �U�����E�    �	�E����E��M�;Ms�U��E��M��������hХ�j�����]����������������������������������������������������������������������������U��EP�MQ�UR�EP�MQ�������]����������������U��EP�MQ�UR�EP�MQ����]�������������������U���0  ���3ŉE��}�t�EP�������ǅ����    jLj ������Q��������������������0���������ǅ����    ǅ����    ������������������������������������f������f������f������f������f������f�������������ǅ0���  �M�������U�������E�H��������U�������E�������M�������  ������������R������������������ u������ u�}�t�EP�������M�3��$�����]����������������������������������������������������������������������������������������U��Q�E�    �X��E��M�Q� �E��E���]����������U��E�X�]����U��Q�X��E��M�Q� �E��}� t�UR�EP�MQ�UR�EP�U�����MQ�UR�EP�MQ�UR������]�������������������������U��j������t�   �)jh �j�������h ��������]����������������������������U��Q�E�    �X��E��M�Q� �E��UR� �E�E�X��E���]���������������������U��j���E�$���E�$�D   ��]����������������U��j���E�$���E�$�   ��]����������������U���8Vh��  h?  �)������E��E%�  =�  t�M���  ���  ��   �U���  ���  u�E����u(�} u"�M���  ���  uE�U����u�} t5�E�P�E�E���$���E�$���E�$�MQj�ۻ����$�b  �U���  ���  t�E%�  =�  u'�M�Q���E�$���E�$�UR�������  h��  �E�P�-������p���  ���]����Au�E���]���]����Au�E���]�E�]����z�E�]���E�]��E��]��E���������Dzh��  �M�Q���������  �E�u��]�E�u��]�E�M�E�M���]ЍU�R���E��$�0�  �$�������E�P���E��$�]�������M��]�u�u����E��$�P������u��}�   ~P�M���   Q���E��$�������]�U�R���E��$���E�$���E�$�EPj�4�����$�   �}����}M�M���   Q���E��$�7������]�U�R���E��$���E�$���E�$�EPj�۹����$�e�M�Q���E��$��������]�U��� th��  �E�P�Y������E��/�-�M�Q���E��$���E�$���E�$�URj�t�����$^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�EP�������]��������������WV�t$�L$�|$�����;�v;��h  �%$�s��  ���   ��  ��3Ʃ   u�%ܪ��  �%$� ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf�����o����   u������r*��$��o��Ǻ   ��r����$��n�$��o��$�o��n�n�n#ъ��F�G�F���G������r���$��o�I #ъ��F���G������r���$��o�#ъ���������r���$��o�I olodo\oToLoDo<o�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��o���o�o�o�o�D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$�$q�����$��p�I �Ǻ   ��r��+��$�(p�$�$q�8p\p�p�F#шG��������r�����$�$q�I �F#шG�F���G������r�����$�$q��F#шG�F�G�F���G�������V�������$�$q�I �p�p�p�p�p qqq�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�$q��4q<qLq`q�D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} u3��  �} t	�E�   ��E�    �E��E��}� u#hܥh�Yj j7h��j��������u̃}� u0�N����    j j7h��h`�hܥ�������   �6  �} t�U;U�  �EPj �MQ��������} t	�E�   ��E�    �U�U��}� u#hx�h�Yj j=h��j�n�������u̃}� u0�����    j j=h��h`�hx��������   �   �M;Mr	�E�   ��E�    �U�U�}� u#h��h�Yj j>h��j��������u̃}� u-�2���� "   j j>h��h`�h���������"   ��   ��MQ�UR�EP������3���]������������������������������������������������������������������������������������������������������������������������̋T$�L$��t�D$�%$�s�L$W�|$��]�T$���   |�%ܪ�����W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$������������������������������������������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+���������������������������������������WV�t$�L$�|$�����;�v;��h  �%$�s��  ���   ��  ��3Ʃ   u�%ܪ��  �%$� ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf����{����   u������r*��$�{��Ǻ   ��r����$�,z�$�({��$��z�<zhz�z#ъ��F�G�F���G������r���$�{�I #ъ��F���G������r���$�{�#ъ���������r���$�{�I {�z�z�z�z�z�z�z�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�{��({0{<{P{�D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$��|�����$�d|�I �Ǻ   ��r��+��$��{�$��|��{�{|�F#шG��������r�����$��|�I �F#шG�F���G������r�����$��|��F#шG�F�G�F���G�������V�������$��|�I h|p|x|�|�|�|�|�|�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��|���|�|�|�|�D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M��EP�M��h����M����E���]� �����������U��Q�M��EP�M��ɦ���M����E���]� �����������U��Q�M��EP�M������M�����E���]� �����������U��Q�M��EP�M��W����M�����E���]� �����������U��Q�M��EP�M��B����M����E���]� �����������U��Q�M��EP�M�������M����E���]� �����������U��Q�M��E�� ̦�M��A    �U��B �E�Q�M�蝢���E���]� ������������������������U��Q�M��E�� ̦�M��U��A�M��A �E���]� ���������������������U��Q�M��E�� ̦�M��A    �U��B �EP�M�蓥���E���]� ��������������������������U��Q�M��E�� ̦�M��A    �U��B �E���]�������������������������U��Q�M��E�� ��M�蕯����]���������������������U��Q�M��E�� ���M�艽����]���������������������U��Q�M��E�� ��M��Y�����]���������������������U��Q�M��E�� ̦�M��`�����]���������������������U��Q�M��E�;Et0�M��1����M�Q��t�E�HQ�M�軠����U��E�H�J�E���]� ������������������������U��Q�M��M�脷���E��t�M�Q�������E���]� ��������������������U��Q�M��M��צ���E��t�M�Q�m������E���]� ��������������������U��Q�M��M�������E��t�M�Q�-������E���]� ��������������������U��Q�M��M������E��t�M�Q��������E���]� ��������������������U����M��} tK�EP���������E��M�Q�������U��B�E��x t�MQ�U�R�E��HQ�������U��B��]� ��������������������������������U��Q�M��E��H��t�U��BP��������M��A    �U��B ��]���������������������������U����M��E��x t�M��Q�U���E�ئ�E���]����������������������U����E������} t	�E�   ��E�    �E�E��}� u#h��h�Yj jYhH�j��������u̃}� u.�T����    j jYhH�hܧh������������   �U�U��E��H��   ta�U�R�*������E��E�P��������M�Q������P��������}	�E������$�U��z tj�E��HQ�������U��B    �E��@    �E���]���������������������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E������} t	�E�   ��E�    �E�E��}� u#h �h�Yj j.hH�j虞������u̃}� u+������    j j.hH�h��h ��7���������W�U�B��@t�M�A    �=�UR�������E�    �EP�	������E��E������   ��MQ�E�����ËE܋M�d�    Y_^[��]���������������������������������������������������������������������������U��Q�} uj �_  ���S�EP���������t����>�M�Q�� @  t.�EP�������P�;�������t	�E�������E�    �E��3���]������������������������������������U����E�    �E�E��M��Q����u|�E��H��  tn�U��E��
+H�M��}� ~Z�U�R�E��HQ�U�R�<�����P�P�����;E�u�E��H��   t�U��B����M��A��U��B�� �M��A�E������U��E��H�
�U��B    �E��]��������������������������������������������������������U��j��   ��]������������������U��j�h �h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} uj �   ���@�EP�������E�    �MQ�֭�����E��E������   ��UR�������ËE�M�d�    Y_^[��]������������������������������������������������������U��j�h �h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    j�������E�    �E�    �	�E���E�M�;����   �U�|��<� ��   �M�|����H��   ��   �U�|���Q�U�R�1������E�   �E�|����B%�   te�}u%�M�|���P聬�������t	�M����M��:�} u4�U�|����Q��t!�E�|���R�C��������u�E������E�    �   ��E�|���R�E�P�������������E������   �j������Ã}u�E����E܋M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������U����E�H���M��U�E��B�}� |�M��%�   �E��M����E���MQ�������E��E���]���������������������������U��j�hP�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E܉E؃}� u#h �h�Yj j)h �j�I�������u̃}� u.�����    j j)h �h`�h ������������  �UR�Y������E�    �E�EԋMԋQ��@��   �E�P�R������E�}��t!�}��t�M����U�����0��U���E���EЊH$�����х�uA�}��t!�}��t�E����M�����0��M���E���ŮB$�� ���ȅ�t	�E�    ��E�   �UȉUă}� u#hp�h�Yj j-h �j��������u̃}� u-�`����    j j-h �h`�hp��������E������}� uP�M�Q���U��E�M��H�}� | �U�����   �M��U����M���UR�M������E��E��E��E������   ��MQ������ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hp�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E܉E؃}� u#h �h�Yj jCh �j�I�������u̃}� u.�����    j jCh �h��h ������������  �UR�Y������E�    �E�EԋMԋQ��@��   �E�P�R������E�}��t!�}��t�M����U�����0��U���E���EЊH$�����х�uA�}��t!�}��t�E����M�����0��M���E���ŮB$�� ���ȅ�t	�E�    ��E�   �UȉUă}� u#hp�h�Yj jGh �j��������u̃}� u-�`����    j jGh �h��hp��������E������}� uP�M�Q���U��E�M��H�}� | �U�����   �M��U����M���UR�M������E��E��E��E������   ��MQ������ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u#h �h�Yj j-h��j�z�������u̃}� u.�����    j j-h��h�h �����������   �} t	�E�   ��E�    �U�U��}� u#h(�h�Yj j.h��j��������u̃}� u+�B����    j j.h��h�h(�����������3�MQ�>������M��Q�U�U�E�M�#Q���t3��������]�������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E܉E؃}� u#h��h�Yj j,hP�j�ɐ������u̃}� u.�
����    j j,hP�h��h���g���������  �UR��������E�    �E�EԋMԋQ��@��   �E�P��������E�}��t!�}��t�M����U�����0��U���E���EЊH$�����х�uA�}��t!�}��t�E����M�����0��M���E���ŮB$�� ���ȅ�t	�E�    ��E�   �UȉUă}� u#hp�h�Yj j0hP�j蟏������u̃}� u-������    j j0hP�h��hp��=������E������}� uZ�M�Q���U��E�M��H�}� |&�U��M��U���   �U��E����U�
��EP�MQ�\������E��U��U��E������   ��EP�"�����ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E܉E؃}� u#h��h�Yj jGhP�j蹍������u̃}� u.������    j jGhP�h��h���W���������  �UR��������E�    �E�EԋMԋQ��@��   �E�P��������E�}��t!�}��t�M����U�����0��U���E���EЊH$�����х�uA�}��t!�}��t�E����M�����0��M���E���ŮB$�� ���ȅ�t	�E�    ��E�   �UȉUă}� u#hp�h�Yj jKhP�j菌������u̃}� u-������    j jKhP�h��hp��-������E������}� uZ�M�Q���U��E�M��H�}� |&�U��M��U���   �U��E����U�
��EP�MQ�L������E��U��U��E������   ��EP������ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u#h �h�Yj j*hЪj�ڊ������u̃}� u.�����    j j*hЪh4�h ��x���������   �} t	�E�   ��E�    �U�U��}� u#h(�h�Yj j+hЪj�a�������u̃}� u+�����    j j+hЪh4�h(������������j �M�QR�P�MQ���������]��������������������������������������������������������������������������������U��j�hЀh�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h �h�Yj j;hH�j�I�������u̃}� u.�����    j j;hH�h��h �������������   �} t�}t�}t	�E�    ��E�   �U܉U؃}� u#hȫh�Yj j<hH�j�Ĉ������u̃}� u+�����    j j<hH�h��hȫ�b���������L�MQ�׾�����E�    �UR�EP�MQ�UR�ؔ�����E��E������   ��EP�{�����ËEԋM�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������U����} u#ht�h�Yj jchH�j薇������u̋M�M��U��B%�   t�} t�}t�}t�����    �����   �M��Q���E��P�}u�M�Q������EU�E�U�E    �U�R�������E��H��   t�U��B����M��A�.�U��B��t#�M��Q��t�E��H��   u
�U��B   �EP�MQ�UR�E�P�*�����P�϶�����E��U�M�#M���u	�E�������E�    �E���]������������������������������������������������������������������������������������U���H�} t�} u3���  �} t	�E�   ��E�    �E�E��}� u#h �h�Yj jqh��j�ׅ������u̃}� u-�����    j jqh��h �h ��u�����3��t  �} t	�E�   ��E�    �U܉U؃}� u#h$�h�Yj jrh��j�_�������u̃}� u-�����    j jrh��h �h$��������3���  ���3��u9Ew	�E�   ��E�    �MԉMЃ}� u#hL�h�Yj jsh��j���������u̃}� u-�!����    j jsh��h �hL��~�����3��}  �E�E�M�M�M��U��U��E�H��  t�U�B�E���E�   �}� �:  �M�Q��  ��   �E�x ��   �M�y }N�U�z }&h��h�Yj h�   h��j��������u̋M�Q�� �E�P�E�+E�3��u��  �M�U�;Qs�E��E��	�M�Q�ŰẺE��M�Q�U�R�E�Q� ������U�+U��U��E�H+M��U�J�E�M��U�
�E�E��E��T  �M�;M���   �U�B%  t �MQ���������t�E�+E�3��u�#  �}� t�E�3��u�E�+E���M��MȋUȉU��E�P�M�Q�UR茶����P蠨�����E�}��u�E�H�� �U�J�E�+E�3��u�   �E�;E�v�M��M���U�UċEĉE��M�+M��M��U�U��U�E�;E�s�M�Q�� �E�P�E�+E�3��u�h�^�M���U��EP�M�Q����������u�E�+E�3��u�;�U���U�E����E��M�y ~�U�B�E���E�   �M��M������E��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t�} u3���   �} t	�E�   ��E�    �E�E��}� u#h �h�Yj jMh��j薀������u̃}� u*������    j jMh��h�h ��4�����3��L�UR誶�����E�    �EP�MQ�UR�EP蜑�����E��E������   ��MQ�N�����ËE܋M�d�    Y_^[��]������������������������������������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E��E܃}� u#h��h�Yj j6hh�j�9������u̃}� u.�z����    j j6hh�ḫh���׽��������/  �}t�} t�}@t	�E�    ��E�   �U؉Uԃ}� u#h�h�Yj j<hh�j�~������u̃}� u.������    j j<hh�ḫh��R���������  �} t
�}@��   �}r�}���w	�E�   ��E�    �MЉM̃}� u#hh�h�Yj j@hh�j�"~������u̃}� u.�c����    j j@hh�ḫhh������������  �E����E�M�M�U�R�#������E�    �E�P�+������M�Q��������U�B%�����M�A�U��t!�E�H���U�J�E���E�E   �b�} uJjxh��j�MQ�{y�����E�} u�\����\��E������J�E�H��  �U�J��E�H��   �U�J�E�M�H�U�E�B�M�U��E��@    �E������   ��M�Q�
�����ËEȋM�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���$�E�E�M�Q��@��   �E�P�O������E��}��t!�}��t�M����U������0��U���E���E��H$�����х�uA�}��t!�}��t�E����M������0��M���E���U�B$�� ���ȅ�t	�E�    ��E�   �U�U�}� u#hp�h�Yj j#h`�j�{������u̃}� u.�]����    j j#h`�h̰hp�躹��������  �M�M��}�t$�U��B��u!�M��Q��   t�E��H��t�����   �U��z u�E�P�V������M��U��;Bu�M��y t����   �U�����M���U��B��@t5�M�����U��E��M���U���M;�t�U�����M������R��U�����E܋M��U܉�E܊M��U��B���M��A�U��B���M��A�U��B���M��A�E%�   ��]��������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h0�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h �h�Yj j/h�j��x������u̃}� u+�
����    j j/h�hP�h ��g���������D�UR�ܮ�����E�    �EP�MQ�˞�����E��E������   ��UR舵����ËE܋M�d�    Y_^[��]������������������������������������������������������������������������������U��Q�=�� u���   ��=��}
���   h�   h�jj���P�������|��=|� u<���   h�   h�jj���Q�������|��=|� u�   �3�E�    �	�U����U��}�}�E���`��M��|�����3���]��������������������������������������������������������U���~��������t�5z��j�|�Q�g������|�    ]����������������������������U��`�]�������U��}`�r?�    k���`�9Mw,�U��`�����R�Mw�����E�H�� �  �U�J��E�� P�  ]�����������������������U��}}#�E��P��v�����M�Q�� �  �E�P��M�� Q�  ]����������������������U��}`�r>�    k���`�9Mw+�U�B%����M�A�U��`�����R�߮������E�� P� ]������������������������U��}}#�E�H������U�J�E��P荮������M�� Q� ]����������������������U����E�E��M�Q�UR�EP�MQ�UR�EP�MQ�N������E��E�    �E���]��������������������������������U����E�E��M�Q�UR�EP�MQ�UR�EP�MQ�������E��E�    �E���]��������������������������������U��E P�MQ�UR�EP�MQ�UR�EP������]������������������������U��j�hP�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t�}t	�E�    ��E�   �E܉E؃}� u#h��h�Yj jth�j�s������u̃}� u.�Թ���    j jth�hx�h���1���������  �} t	�E�   ��E�    �UԉUЃ}� u#h��h�Yj juh�j�s������u̃}� u.�[����    j juh�hx�h��踱��������  j��s�����E�    �$��M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���M̋U�ẺB�M̉M��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H�$�j�U�R�΀�����<3�u&hزh�Yj h�   h�j�r������u��E������G����    ��   �}� tu�U�B���EȋM�UȉQ�EȉE��M�;$�tM�U�z t�E�H�U���M��E�H�J�U��    �E�$��H�$��E��M�$��h�   hD�jj�{m�����E�}� u�E�����薷���    �L�U��    �E�$��H�=$� t�$��E��M��A   �E�   �U�E�B�M�$��E������   �j�0�����ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��\"  迼�����3ŉE�ǅ����    ǅ����    ǅ����    �} u
�   �S  ������P�MQj�, ��u
ǅ����    �   i�  ������������
  s��7���3ɋ�����f������h  ������P������Q�( ��u8j h_  h�ht�h��h$�h  ������R�5�����P��y����������������������Q蝘������@vo������R艘�����������TA�������j hh  h�ht�h`�j�`�P������������+����  +���P������Q�xz����P�Cy�����} t*�UR��������@v�EP�������M�TA�������莴��� ������聴���     �}uǅ����p��
ǅ�������   k� �E���t�U�������
ǅ�������   k� �U�
��t�}uǅ�������
ǅ�������   k� �E���tǅ�������
ǅ�������} t�U�������
ǅ�������} tǅ�������
ǅ�������} t�E�������
ǅ�������} tǅ�������
ǅ������������ t�������������'�} t�U�������
ǅ������������������������ tǅ����|��
ǅ�������} tǅ����Զ�
ǅ������������Q������R������P������Q������R������P������Q������R������P������Q������R������P�M�� �Rh�h�  h   ������P�������D������������ }*j h  h�ht�h��j"j�M����Q�fi���� �=���������������� }8j h�  h�ht�h�h��h   ������P�ײ����P�tv����h  h �������Q�#�����������������uj�vy����j�nm��������u�   �3��M�3�������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��} u��EP�MQ�UR�EP�MQ�<���]�����������U��} t�E;Et�M;Mt�E��U$R�E P�MQ�UR�EP������E]���������������������U��Q�M��E��@ �} ��   �ϛ���M��A�U��B�M��Pl��E��H�U��Ah�B�M��;4�t�E��H�Qp# �u
�0����M���U��B;|�t�M��Q�Bp# �u�O����M��A�U��B�Hp��u�U��B�Hp���U��B�Hp�M��A��U��J�U���J�E���]� ���������������������������������������������������������U��Q�M��E��H��t�U��B�Hp����U��B�Hp��]����������������������U��Q�M��E���]�������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j��h�����E�    h��h�_j j j j �,h������u̃} t�M��U�|��E���M��U�}� �0  �E�;E��$  �M�Q����  ��t)�E�H����  t�U�B%��  ��u�l���u��  �U�z tyj j�E�HQ�Q�������tj�U�BP��  ����t$�M�QRh��j j j j �`g������u��)�M�QR�E�HQh��j j j j �5g������u̋E�HQh��j j j j �g������u̋E�H����  ����   �U�BP�M�Q������  R�E�� Ph��j j j j ��f���� ��u̃=h� t3�U�BP�M�� Q��  ����u�U�BP�M�� Q�h�����U�R�EP�7  ���   �M�yu;�U�BP�M�� Qh8�j j j j �Bf������u̋E�P�MQ�A7  ���Y�U�B%��  ��uI�M�QR�E�H������  Q�U�� Rhh�j j j j ��e���� ��u̋M�Q�UR��6  �������E������   �j譞�����h��h�_j j j j �e������u̋M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hЂh�Ld�    P���SVW���1E�3�P�E�d�    �e��E�    3��E��E��E��E��EĉEȉẺEЍM�Q�4 �U��U؃} ��   �} u
�   �   �E�E��M�U��D
��E܋M�;M�s	�   �v�r�E�    �U���E�M؃���#M��M��U؃���#U܉U܋E�;E�t�M�M؉M��U���E����E������#�   Ëe��E�   �E������E��	�E�����3��M�d�    Y_^[��]�����������������������������������������������������������������������������������������U����E�E��M���M�}� t'�U��E��M�M�U���U�E�;E�t3���ĸ   ��]����������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�   �l���u
�   ��  j�c�����E�    �Q����Eԃ}����   �}����   �MԉM܋U܃��U܃}���   �E��$�T�h�h�_j j j j �)b������u��   h4�h�_j j j j �b������u��dh`�h�_j j j j ��a������u��Bh��h�_j j j j ��a������u�� h��h�_j j j j �a������u��E�    ��  �|��E���M��U�}� ��  �E�   �E�H����  ��t#�U�zt�E�H����  ��t	�U�zu�E�H����  ��X��U���E���j�t�P�M��Q���������uz�U�z t=�E�HQ�U�BP�M�� Q�U�BP�M�Qhȿj j j j �`����(��u��-�E�� P�M�QR�E�Ph��j j j j �`���� ��u��E�    j�t�R�E�H�U�D
 P�$�������uz�M�y t=�U�BP�M�QR�E�� P�M�QR�E�Ph@�j j j j �`����(��u��-�U�� R�E�HQ�U�Rh�j j j j ��_���� ��u��E�    �M�y ��   �U�BP�v�Q�U�� R�{�������ud�E�x t2�M�QR�E�HQ�U�� Rh��j j j j �_���� ��u��"�M�� Qh��j j j j �[_������u��E�    �}� uz�E�x t=�M�QR�E�HQ�U�BP�M�� Q�U�RhP�j j j j �
_����(��u��-�M�QR�E�� P�M�Qh��j j j j ��^���� ��u��E�    �G����E������   �j誗����ËEЋM�d�    Y_^[��]Ð���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h0�h�Ld�    P���SVW���1E�3�P�E�d�    �} t	�E�   ��E�    �E��E܃}� u&h��h�Yj h�  h��j�\������u̃}� u+�ޢ���    j h�  h��h��h���8������s�l���u�fj�D]�����E�    �|��E���M��U�}� t$�E�H����  ��u�UR�E�� P�U�����E������   �j�L�����ËM�d�    Y_^[��]�����������������������������������������������������������������������������������U���8���3ŉE��E�P�}������   ���|� u'�   �� �|� u�l���t?�   ��|� t1h��h�_j j j j �[������u�j 躚�����   �3��M�3���y����]����������������������������������������������U��h�]�������U��`�]�������U��h�]�������U��j�hP�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�     �} t	�M�    �} t	�U�    �EP贂������u3���   j�[�����E�    �M�� �M�U�B%��  ��t"�M�yt�U�B%��  ��t	�M�yukj�UR�EP�ډ������tU�M�Q;UuJ�E�H;p�<�} t�U�E�H�
�} t�U�E�H�
�} t�U�E�H�
�E�   ��E�    �E������   �j蟒����ËE��M�d�    Y_^[��]���������������������������������������������������������������������������������������������������U��} u3��1j j �E�� P�ʈ������u3���M�� Qj ���R�0 ]�����������������U��Q�} t	�E�   ��E�    �E���]����������������U��j�hp�h�Ld�    P���SVW���1E�3�P�E�d�    �} t	�E�   ��E�    �E܉E؃}� u&h$�h�Yj h�  h��j��W������u̃}� u.�����    j h�  h��hH�h$��x������m  j�X�����E�    �U�|���E�    �	�M����M��}�}�U��E�D�    �M��U�D�    �ӡ|��E���M��U�}� ��   �E�H����  |f�U�B%��  ��}V�M�Q����  �E�L����U�B%��  �U�L��E�H����  �U�D��M�A�U�J����  �U�D��W�E�x t/�M�QR�E�HQ�U�Rht�j j j j ��V���� ��u���M�Qh��j j j j ��V������u������E�x��H,�U�p��B0�E������   �j菏����ËM�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������U��� V�E�    �} t	�E�   ��E�    �E��E�}� u&h$�h�Yj h�  h��j�?U������u̃}� u0耛���    j h�  h��h��h$��ړ����3���  �} t	�E�   ��E�    �U��U�}� u&h�h�Yj h�  h��j��T������u̃}� u0�����    j h�  h��h��h��\�����3��E  �} t	�E�   ��E�    �M�M�}� u&h<�h�Yj h�  h��j�CT������u̃}� u0脚���    j h�  h��h��h<��ޒ����3���   �E�    �	�E����E��}�}�M��U�E��u�L�+L��U��E�L��M��U�E��u�L�+L��U��E�L��M��U�|� u�E��M�|� t$�}� t�}�u�}�u�l���t�E�   �r����E�M�P,+Q,�E�P,�M�U�A0+B0�M�A0�U�    �E�^��]�������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    �E�P�M��L\���M�蒟��P�MQ�E������M��yl����]�����������������������U����} t	�E�   ��E�    �E��E�}� u&h$�h�Yj h
  h��j�R������u̃}� u.�H����    j h
  h��h��h$�袐�����   �E�    �	�U����U��}�}>�E���X�Q�U��E�L�Q�U��E�L�Qh�j j j j ��Q���� ��u�볋E�H,Qh4�j j j j �Q������u̋E�H0Qh\�j j j j �Q������u̋�]���������������������������������������������������������������������������������U��Q�EP�[y������u�����M�� �M��U��B��]���������������������U��Q�h��E��M�h��E���]���������������������U��Q�d��E��M�d��E���]���������������������U��Q�`��E��E���]��������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    j��P�����E�    �EP�^x������tj�M�� �M�U�B%��  ��tH�M�yt?�U�B%��  ��t/�M�yt&hh�h�Yj h?  h��j�sO������u̋E�M�H�E������   �j褈����ËM�d�    Y_^[��]�����������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �l��E܃}�t�M����  ���t	�E�    ��E�   �U�U��}� u&h��h�Yj hw  h��j�wN������u̃}� u0踔���    j hw  h��h��h���������l��sj�&O�����E�    �l��M܃}�t7�U��t�d�   ��E��%��  �d��l�    �M�l��E������   �j�$�����ËE܋M�d�    Y_^[��]����������������������������������������������������������������������������������������U��Q�h��E��M�h��E���]���������������������U��Q�h��E��M�h��E���]���������������������U��EP��f����]����������������U��Q�} u�   �E������E�j�t�Q�U��R���������t!�EPh �j j j j��L������u��Lj�u�R�E���P��������u�MQh��j j j j�L������u�j�E��Q��Z������]��������������������������������������������������������U��j j j �EP�MQ�L����]����������������������U��EP�MQj �UR�EP�\L����]������������������U��EP�MQ�UR������]��������U���$�E�    �E�    �E�    �E�    �E�    �} t	�E�   ��E�    �E�E��}� u&ht�h�Yj h  h��j�K������u̃}� u.�U����    j h  h��h��ht�诉��������w�E�    �U������U��E��Q�PT�����E�U��E+�E�3�+M���M�}v�U�U���E�   �E���E�M�U�D
+E��E��M�+M�+M��M܋E܋�]���������������������������������������������������������������������������������U��j j �EP�MQ�UR�J����]��������������������U���,�E��#Eu	�E�   ��E�    �M��M�}� u&h��h�Yj h@  h��j�I������u̃}� u0�ӏ���    j h@  h��h��h���-�����3��E  �} t�E;Er	�E�    ��E�   �M��M�}� u&h��h�Yj hA  h��j�I������u̃}� u0�M����    j hA  h��h��h��觇����3��   �}v�E�E���E�   �M���M3�+U���U܋E�M܍T�U��EE��E�M;M�v�֎���    3��i�UR�EPj�M�Q�D�����E��}� u3��F�U�U�U�E��#�+U�UԋM�+M܃��M�j�u�R�E؃�P�1o�����M؋U���Eԋ�]�������������������������������������������������������������������������������������������������������������������������������U��j j �EP�MQ�UR�EP�'�����]����������������U���8�} u!�EP�MQ�UR�EP�MQ��G������  �} u�UR�a����3��  �E������E�j�t�Q�U��R��������t1�EPh8�j j j j�6G������u������    3��_  j�u�R�E���P���������u�MQh��j j j j��F������u̋E��#Eu	�E�   ��E�    �M��M�}� u&h��h�Yj h�  h��j�<F������u̃}� u0�}����    j h�  h��h��h���ׄ����3��  �} t�E;Er	�E�    ��E�   �M�M�}� u&h��h�Yj h�  h��j�E������u̃}� u0������    j h�  h��h��h���Q�����3��  �E��Q�O�����U��M+
+��Ẽ}v�U�U���E�   �E����E3�+M���MԋU�EԍL�M؋UU؉U܋E;E�v�e����    3��   �MQ�URj�E�P�A�����E��}� u3��   �M�M�M�U��#�+M�M�E�+Eԃ��E�j�u�Q�UЃ�R�k�����EЋM���U�;Uv�E�E���M̉MȋU�R�EP�M�Q�M����j�U��P�S�����E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j j �EP�MQ�UR�EP�MQ�7K����]������������U����E�    �E�    �E�    �} v�����3��u;Es�|����    3��s�E�E�E��} t�MQ�UR�EP�a������E��M Q�UR�EP�MQ�U�R�EP萐�����E�}� t �M�;M�s�U�+U�Rj �E�E�P��i�����E��]�����������������������������������������������������������U��j j j �EP�MQ�UR�	�����]������������������U��EP�MQj �UR�EP�MQ�Տ����]��������������U��j j j �EP�MQ�UR�EP�I����]��������������U��EP�MQj �UR�EP�MQ�UR�I����]����������U����E�    �E�P�MQ�UR�EP�MQ�UR��i�����E��}� u�}� t�������t
跇���M���E���]���������������������������U��Q�} v�����3��u;Es�s����    3��K�E�E�E�MQ�UR�EP�MQ���R�EP��  ���E��}� t�MQj �U�R��g�����E���]������������������������������������������U��Qj j j�EP�MQ��U�����E��E���]�������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E��E܃}� u&h��h�Yj h�  h��j��?������u̃}� u-�7����    j h�  h��hоh���~����3��c�}�v�����    3��Nj�@�����E�    j �UR�EP�MQ�UR�EP��  ���E��E������   �j�x����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������U��j�h��h�Ld�    P��SVW���1E�3�P�E�d�    j�?�����E�    �EP�MQ��p�����E������   �j��w����ËM�d�    Y_^[��]�������������������������������������U��Q�=d� vZ�d���9l�u;�u]����u&h��h�Yj h  h��j�>������u��l�    ��l����l��} u�  �}uOj�u�P�M�����Q���������t/�URh�j j j j�>������u�������    �5  �=h� tDj j j �MQj �URj�h�����u%hH�h�_j j j j �=������u���  �MQ��e������u&hp�h�Yj h*  h��j�=������u̋E�� �E��M��Q����  ��tI�E��xt@�M��Q����  ��t/�E��xt&hh�h�Yj h0  h��j�<������u̋l����m  j�t�P�M���Q����������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��X�Phȿj j j j�<����(��u��<�U��� R�E��HQ�U��B%��  ��X�Qh��j j j j�U<���� ��u�j�t�P�M��Q�E��L Q�����������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��X�Ph@�j j j j��;����(��u��<�U��� R�E��HQ�U��B%��  ��X�Qh�j j j j�;���� ��u̋E��xuj�M��y����u	�U��z t&h��h�Yj hi  h��j��:������u̋M��Q��$R�v�P�M�Q��a�����U�R�vs�����`  �E��xu�}u�E   �M��Q;Ut&h<�h�Yj hw  h��j�:������u̋M��t�+Q�t��l�����   �M��9 t�U���M��Q�P�;���;E�t&h��h�Yj h�  h��j�:������u̋U��B����M��y t�U��B�M����:�|�;E�t&h��h�Yj h�  h��j��9������u̋U���|��M��Q��$R�v�P�M�Q�`�����U�R�;r�����(�E��@    �M��QR�v�P�M��� Q�x`������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�EP�Ej����]��������������U��j j j�EP��l����]����������U����E�    �E�P�MQ�UR�EP�MQ�J   ���E��}� u�}� t��}����t
��}���U���E���]�������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    j�8�����E�    �=d� vZ�d���9l�u;�:V����u&h��h�Yj h  h��j��6������u��l�    ��l����l��p��E��=d��t�M�;d�u̃=h� tu�UR�EP�M�Q�UR�EPj j�h�����uP�} t%�MQ�URh �j j j j �6������u�� h`�h�_j j j j �6������u��D  �U����  ��t�l���u�E�   �}�v3�MQh��j j j j�C6������u̃} t	�E�    ��  �M����  ��t:�}t4�U����  ��t&�}t h��h�_j j j j��5������u̋M��$�MԋU�R�S�����E�}� u�} t	�E�    �r  �p����p��}� tI�U��    �E��@    �M��A    �U��B�����E�M�H�U��B   �E��@    �   ���+p�;Mv�p�U�p��
�p������t�E�t��t�;x�v�t��x��=|� t�|��M�H�	�U����E�|���U��B    �E�M�H�U�E�B�M�U�Q�E�M�H�U�E��B�M�|�j�t�R�E��P�4[����j�t�Q�U�E�L Q�[�����UR�w�P�M�� Q��Z�����U�� �U��E������   �j�m����ËE؋M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�EP�MQ�UR���P�MQ�m�����E��E���]���������������������U��j�EP�_����]��������������U��j�hЁh�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E��E܃}� u&h��h�Yj h�  h��j��1������u̃}� u1�'x���    j h�  h��h��h���p��������G  �=d� v[�d���9l�u;��P����u&h��h�Yj h�  h��j�f1������u��l�    ��l����l�j�02�����E�    �UR�Y������u&hp�h�Yj h�  h��j�1������u̋M�� �M�U�B%��  ��tH�M�yt?�U�B%��  ��t/�M�yt&hh�h�Yj h�  h��j�0������u̋E�xu�}u�E   �M�Q�U��E������   �j�i����ËE؋M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������U��j j j�EP�MQ�j����]����������������������U����E�    �E�P�MQ�UR�EP�MQ�UR�F   ���E��}� u�}� t�u����t
�u���M���E���]���������������������������U��Q�EP�MQ�UR�EP�MQ�������E��}� t�E��?�} u�} t	�U�   �E��%�EP�Qg������u�} t	�M�   3��뗋�]��������������������������������U���x���3ŉE��EP�M��98���E�    �	�M����M��U�z}�E�H�M���E�   �U�;U���   �EE��H �M��M��:{����t0�M��.{����zt~ �M��{��PhW  �E�P�B�����E��hW  �M�Q�M���z��P��)�����E��}� t	�U��U���E�    �E��M��L��t����U���s���     �E�Phd�kM��1   +�RkE��L�Q�g������}*j h	  h��hl�h��j"j�s���R��*���� �s���M��������U��U��}�s���k���E��D� �M�Q�U�Rh��j j j j �b-������u̍M��G���M�3��K����]�������������������������������������������������������������������������������������������������������������������������U��j�hp�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j�#-�����E�    j�EP�MQ�UR�EP�MQ�}  ���E��E������   �j�Fe����ËE�M�d�    Y_^[��]������������������������������������������U��Qj j j�EP�MQ�UR�Ns�����E��E���]�������������������������U����E�    �E�    �E�    �} v�����3��u;Es�q���    3��g�E�E�E��} t�MQ�4�����E��UR�EP�MQ�U�R�EP��?�����E�}� t �M�;M�s�U�+U�Rj �E�E�P��Q�����E��]�������������������������������������������������������U����E�    �E��M��} u�UR�EP�MQ�U�R�~&������  �} t�}� u�EP�MQ��8����3��  �=d� v[�d���9l�u;�MI����u&h��h�Yj h�  h��j��)������u��l�    ��l����l��p��U�=d��t�E�;d�u̃=h� ty�MQ�UR�E�P�MQ�U�R�EPj�h�����uR�} t%�MQ�URh�j j j j �)������u�� h4�h�_j j j j �)������u�3��  �}��v`�} t)�UR�EP�M�Qh`�j j j j�b)���� ��u���E�Ph��j j j j�A)������u��)o���    3��A  �}th�U����  ��tZ�E%��  ��tM�} t%�MQ�URh��j j j j��(������u�� h��h�_j j j j��(������u��Qj�u�R�E�����P�d�������t1�MQh�j j j j�(������u��jn���    3��  �EP�P������u&hp�h�Yj h  h��j��'������u̋U�� �U�E�xu�E�   �}� t=�M�y����u	�U�z t&hȼh�Yj h#  h��j�'������u��d�M�Q����  ��u�E%��  ��u�E   �M�p�;Qs1�EPhp�j j j j�'������u��tm���    3��  �} t%�U���$R�E�P��u�����E��}� u3��c  �#�M���$Q�U�R�H�����E��}� u3��>  �p����p��}� u{�=p��s;�M��p�+Q�p����+p�;E�v�p�M��p��
�p������U��t�+B�t��t�M��t��t�;x�v
�t��x��M��� �M�U��E�;Bv$�M��U�+QR�w�P�M��U�QR�M����j�t�P�M�M�Q��L�����}� u�U��E�B�M��U�Q�E��M�H�U��E��B�} u4�} u�M�;M�t&h��h�Yj h�  h��j�%������u̋E�;E�t�}� t�E���   �M��9 t�U���M��Q�P�;���;E�t&h(�h�Yj h�  h��j�,%������u̋U��B����M��y t�U��B�M����:�|�;E�t&hd�h�Yj h�  h��j��$������u̋U���|��=|� t�|��U��Q��E�����M��|���E��@    �M��|��E��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;��u����K�������������������U���,VW�   ����}��E�E��}� t:�M����t0�E��M��U����U��E��E�M��B�E��M�Q�U��H �ыU�U�E��E��}� t�M����t�E� @��E�P�M�Q�U�R�E�P�8 _^��]� ��������������������������������������������������U��Q��E�H3M��@��j �MQ�U�BP�M�QRj �EP�M�QR�EP��a���� �E��E���]�����������������������U��QS��E�H3M�e@���M�Q��ft�E�@$   �   �v�tj�M�QR�E�HQ�U�BPj �MQ�U�BP�MQ�?a���� �U�z$ u�EP�MQ�?a��j j j j j �U�Rh#  �#�����E��]�c�k ��   [��]������������������������������������������������������U����E�    �E�����M�3��E�U�U��E�E�M���M�d�    �E�E�d�    �UR�EP�MQ�o���E��E�d�    �E���]�������������������������������������XY�$�����������XY�$�����������XY�$�����������U���8S�}#  u�<�M��   ��   �E�    �E������M�3��EЋU�UԋE�E؋M�M܋U �U��E�    �E�    �E�    �e�m�d�    �EȍE�d�    �E�   �E�E��M�M���Q�����   �U��E�P�M�R�U����E�    �}� td�    ��]ȉd�    �	�E�d�    �E�[��]�����������������������������������������������������������������������U����MSVW�q�ދ}�A�E��u���x>�M���u�+j���M�U�N��9L��U�}�U�;L��U�~���uO�u��څ�yȋM�EF�0�E�;Yw;�v��i���M���_^[����]�����������������������������������������U��QS�E���E�d�    �d�    �E�]�m��c���[��]� ��������������U���SVWd�5    �u��E��j �EP�M�Q�UR�< �E�H����U�Jd�=    �]��;d�    _^[��]� �����������������������U��MV�u��O�����   �N�O�����   ��^]�����������������������U��V�O���u;��   u�sO���N^���   ]��bO�����   �y t�A;�t�ȃy u�^]�mh���F�A^]����������������������������U���O�����   ��t�M9t�@��u��   ]�3�]����������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�R\���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�\���� �E�_^[�E���]���������������������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�[���� �E�_^[�E���]���������������������U��E�HQ�   k� �M�T(Rj �E�HQ�����]� ����������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ����������������������������U��Q�M��E�� ���E���]� �������U��Q�M��E�� ���M�Q��C������]�����������������U��Q�M��E���]� ����������������U����M��E���	P�M��	Q��D������t	�E�    ��E�   �E���]� ��������������������U����M��E���	P�M��	Q�D������t	�E�   ��E�    �E���]� ��������������������U��Q�M��M������E��t�M�Q�=h�����E���]� ��������������������U��Q�M��EP�M�Q��F������]� �������������������U��Q�M��E�P��Y������]����������U����M��E���	P�M��	Q��C������~	�E�   ��E�    �E���]� ��������������������U��Q�M��EP�M�Q�E"������]� �������������������U��Q�M��E�����]����������������U���!M���} t��`����]����������U��Q����E��M����E���]���������������������U��   k� ǁ0��S�   �� ǂ0��N�   ��ǀ0�
k�   k�ǂ0�4_�   ��ǀ0��[�   k�ǂ0��S�   k�ǁ0��C�   k�ǀ0��j�   ��ǁ0��L�   k�	ǀ0�T:]���������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �}��   �����u3���  �u ����u�	��3���  ��&���@ �(��a2������P����}�cJ������3��  �Z3����|�J0����|j ��/������t�^F���-J�����3��g  j�,�������������F  �} ��   �=�� ~{���������E�    �=�� u�<��� 4��j���;������ tj �������N����E���I������E������   ��} u�=|��t�zI����3��   �   �}��   �|�R��.�����E�}� uxh�   h�jh�  j�G.�����E�}� tP�E�P�|�Q�������t%j �U�R��+�����D �M��U��B�����j�E�P�!$����3���3����}u
j �d�����   �M�d�    Y_^[��]� ������������������������������������������������������������������������������������������������������������������������������������������������������������U��}u�9���EP�MQ�UR�   ��]� ����������U��j�h0�h�Ld�    P���SVW���1E�3�P�E�d�    �e��E�   �} u�=�� u3��Z  �E�    �}t�}uT�=� t�EP�MQ�UR���E�}� t�EP�MQ�UR�,���E�}� u�E�    �E������E���   �EP�MQ�UR�6���E�}u=�}� u7�EPj �MQ��5���URj �EP�-,���=� t�MQj �UR���} t�}u@�EP�MQ�UR��+����u�E�    �}� t�=� t�EP�MQ�UR���E��E������D�E���U܋E�P�M�Q�UR�EP�MQ��a����Ëe��E�    �E������E��
�E������E�M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������U��}u�EPj �MQ��*���UR�EP�\����]�����������������������U��Qj j j���P�MQ��L�����E��E���]�����������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_������������������������������������������������������������������������̀�@s�� s����Ë���������������������������̹   �-x���   �-����   �-x�f~�%���=  ��L  �Z���u���f/�v
�   �=  f/��!  �5p�f/��  fo�fs�fs���t:���f/�w,fW�f/�t"P��<$f�$f� Xu�   ��   3��   ��fW�f/���   �P��%X�fn-��fo���� fo�f��f��fs�4fo�f��fo�f��fo�f��fo�f��ff�fb�f��f��f��f��f��f��f��f��f~��� ~#f��f��f~�fs�f~��t
�   �    f~�fs�f~�ú   �   3��   �Ã� ��<$�$��t����u(�-���$�D$    �D$�D$�D$����؃� ù   �-x���   �-����   �-x�fo�fs�f~�%���=  ��b���������fo�fs�fs����f/�v/��t�   �@����   �6�����   �*����   � ������f/�s'fW�f/��0����   ������   ���������fo؃�u�x�f/�rf\�fo�fs�#fs�#f~��t
�   ����f/�������p�f/������������u�*�����@��X��fn%��fn-��fn5��fn�fn�fb��    ��+�fn�f��fo�fs�3fs�3fo�fs�fs�ff�fb�f��ff�fb�f��f��fs�4f��Ë���;�u�*�Å��Y����=`��ك� ���E���V�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U������]�h��  h?  �;�����E��E%�  =�  ��   ���E�$�I6�����E��}�t�}�t!�}�t3�Jh��  �M�Q�5;�����E�   h��  �U�R�;�����E���i�E�P���E�$j�i4�����P�M�Q�E��`���$���E�$jj�
�����&�U������U�E�E�h��  �M�Q�:�����E���]����������������������������������������������������������������������̃��$� ���   ��ÍT$���R��<$�D$tQf�<$t��L���   �u���=�� �����   ����<H���  �u,��� u%�|$ u���:���"��� u�|$ u�%   �t����-�|�   �=�� �d���   ������Z�������������������������������������������������������U��E�<Ű� u�MQ�'T������u
j������U�հ�P�  ]��������������������U�������u�EPj �H h�   ��2����]����������U����E�    �	�E����E��}�$}O�M��<Ͱ� t@�U��<մ�t3�E��Ű��M��U�R� j�E�P�C�����M��Ͱ�    ��E�    �	�U����U��}�$}3�E��<Ű� t$�M��<ʹ�u�U��հ��E�M�Q� 뾋�]�����������������������������������������������������U��j�hP�h�Ld�    P���SVW���1E�3�P�E�d�    �E�   �=�� u�G��j�1����h�   �1�����E�<Ű� t
�   �   h  h��jj������E�}� u��M���    3��jj
�Y�����E�    �M�<Ͱ� u"j h�  �U�R��5�����E�M�Ű��j�U�R�������E������   �j
�`@����ËE��M�d�    Y_^[��]������������������������������������������������������������������������������������U����E�    �E�    �	�E����E��}�$}F�M��<ʹ�u7kU�� ��E��Ű��M����M�j h�  �U��հ�P��4����뫸   ��]���������������������������������������������U��E�Ű�Q� ]�����������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �e�} t8�E�8csm�u-�M�yu$�U�z �t�E�x!�t�M�y"�t�   �U�z ��   �E�H�y tS�E�    �U�B�HQ�U�BP�+���E������+�M��t	�E�   ��E�    �E�Ëe������E������,�U�B���t�U�B��M�}� t�U��M�Q�P�ҋM�d�    Y_^[��]���������������������������������������������������������������������������������U��Q�M��EP�M��G���M����E���]� �����������U��Q�M��EP�M��W���M����E���]� �����������U��Q�M��E�� ��M��9����]���������������������U��Q�M��M�����E��t�M�Q�R�����E���]� ��������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �e�E�E��E�    �   k���E��M̋U�BP�M�Q�	�����E��5�����   �U��r5�����   �E��d5���M���   �V5���U���   �E�    �E�   �E�   �E P�MQ�UR�EP�MQ�C�����E��E�    ��   �U�R�  ��Ëe���4��ǀ�      �E�H�MЋU�z�   �E�H���   �щU��	�E�H�MԋUԉU��E�H�M��E�    �	�U���U�E�M�;HsAkU��E؋M�;L~/kU��E؋M�;LkU��E؋L���M��U��EЋЉM��뫋U�R�EPj �MQ������E�    �E�    �E������E�    �   �   �   k���M�Ủ�E�P��������3���Mĉ��   ��3���U����   �E�8csm�u\�M�yuS�U�z �t�E�x!�t�M�y"�u/�}� u)�}� t#�U�BP�6������t�M�Q�UR�����ËE܋M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h d�    PQSVW���3�P�E�d�    �e��~2�����    u��K���E�    ����]2���M���   j j �3����%��E�������E���������M�d�    Y_^[��]���������������������������������������������������U����E�E��}  t�M Q�UR�E�P�MQ�BF�����}, u�UR�EP�j?����MQ�U,R�[?���E$�Q�UR�EP�M�Q�Z�����U$�B���M�Ah   �U(R�E�HQ�UR�EP�M�Q�UR�f������E��}� t�EP�M�Q������]����������������������������������������������������������U��Q�E��M��U��:csm�uN�E��xuE�M��y �t�U��z!�t�E��x"�u!�M��y u�0��ǀ�     �   ��3���]��������������������������������������U���D�E� �E� �E�x�   �M�Q���   �E��	�M�Q�U܋E܉E�}��|�M�U�;Q}��DI���E�8csm��[  �M�y�N  �U�z �t�E�x!�t�M�y"��&  �U�z �  ��/�����    u�  �/�����   �E�/�����   �M�E�j�UR�$������t��H���E�8csm�u;�M�yu2�U�z �t�E�x!�t�M�y"�u�U�z u�aH���//�����    ty�!/�����   �E��/��ǀ�       �M�Q�UR�  ������t�C�M�Q�K  ���Ѕ�t+j�EP������h$��M��v��h���M�Q�w/����.����U�:csm���  �E�x��  �M�y �t�U�z!�t�E�x"��i  �M�y �5  �U�R�E�P�M�Q�U R�EP�8�����E���M���M�U����U��E�;E���   �M��;U��E��M�;H~�˺   k� �M�A�E��U��B�E���M���M�U����U��}� ��   �E�H�Q���U��E�H�Q��E���M���M�U����U��}� ~d�E���MԋU�BP�M�Q�U�R�f������u���E��E�P�M$Q�U R�E�P�M�Q�U�R�EP�MQ�UR�EP�MQ�P�����,�	���D���������(�U�%���=!�r��<F���M�y t��,F���U��tj�EP������M�����   �U�%���=!���   �M�y ��   �U�BP�MQ�/  ���Ѕ���   �,�����   �E��,�����   �M��|,���U���   �n,���M���   �}$ u�UR�EP�:����MQ�U$R��9��j��EP�MQ�UR�������E�HQ�u������,���U���   �,���M���   �@�U�z v7�E��u*�M$Q�U R�E�P�MQ�UR�EP�MQ�UR�^  �� ��A����+�����    u���D����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���V�E�8  �u�o  �P*�����    tZ�B*����j � 9��   tC�M�9MOC�t8�U�:RCC�t-�E$P�M Q�UR�EP�MQ�UR�EP��������t�  �M�y t��
C���U�R�E�P�MQ�U R�EP�3�����E���M����M��U����U��E�;E���   �M��U;|e�E��M;HZ�U��B�����M��Q�| t'�E��H�����U��B�L�   k� �L��u�U��B�����M��Q���@t�n���j�M$Q�U R�E�Pj �M��Q�����E�PR�MQ�UR�EP�MQ�UR������,�*���^��]������������������������������������������������������������������������������������������������������U����} t��A���} u������E� �E�    �	�E����E��M�U�;}m�E�H�Q���U��E�H�Q��E���M���M�U����U��}� ~4�E���M�U�BP�M�Q�U����EPR��������t�E���뀊E���]�����������������������������������������������U��Q�E�    �	�E����E��M�U�;}'h���E����M�Q�L� ������t����2���]��������������������U��Q�3'�����    t	�E�   ��E�    �E���]������������������������U����} t��@���E��M��}� t��@���U��:csm�u/�E��xu&�M��y �t�U��z!�t�E��x"�u���?���M��Q�B���E�M��Q�B��M���U����U��E���E�}� ~0�M��U��E��H��Q�M����P�i������u�   ��3���]�������������������������������������������������������������U��E�P�]����U��Q�E�M�M��U�z |'�E�H�U�
�M�Q�M��M��U�E�B�E��E���]���������������������������U��j�hЃh�Ld�    P���SVW���1E�3�P�E�d�    �e�E���   �t�U�U���E�H�U�D
�E��E�    �MQ�UR�EP�MQ�s2�����E��}�t�}�t+�R�U��R�E�HQ�_����P�U�BP�M�Q�4����)j�U��R�E�HQ�4����P�U�BP�M�Q�V>���E�������   Ëe������E������M�d�    Y_^[��]�����������������������������������������������������������������������U��j�hp�h�Ld�    P���SVW���1E�3�P�E�d�    �e��E�    �E�x t-�M�Q�   k� �T
��t�E�x u�M���   �u3��j  �E���   �t�U�U���E�H�U�D
�E��E�    �M���   tn�E���td�=P� t[�P��E�j�U�R�`������t6j�E�P�J������t$�M�U܉�E��P�M�R������M���@<���  �U���tXj�M�QR�������t9j�E�P��������t'�M�U�B��M��Q�U�P�>�����M����;���@  �U���txj�M�QR�������tYj�E�P�������tG�M�QR�E�HQ�U�R�������E�xu"�M�9 t�U��R�E�Q������U���\;���   �E�x uZj�M�QR�������t>j�E�P�������t,�M�QR�E��P�M�QR�^����P�E�P���������:���[j�M�QR��������tAj�E�P�������t/�M�QR�.������t�E���t	�E�   ��E�   ��:���E�������   Ëe�������E������E��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} u3��l�E��M��U��:csm�uW�E��xuN�M��y �t�U��z!�t�E��x"�u*�M��y u!� ���   �E��U�����M���   �3���]���������������������������������U���(�} u3���  �E��M��} t�   k� �M�T����   �E��8MOC�t�M��9RCC�t�U��@uz�E��8csm�uK�M��yuB�U��z �t�E��x!�t�M��y"�u�U��z u�?�����    u3��H  �*���   �E��E�����U��
�   �$  �E��8csm��  �M��y�  �U��z �t�E��x!�t�M��y"���   �U��z u#������    u3���   ������   �E��M�M܋U�U؋E�   ��E؋M��Q�B���E�M��Q�B��M���U����U��E���E�}� ~d�M��U�E��HQ�U�R�E�P��������t?�%���   �E�M����E��} t�M�Q�U�R�EP�M�Q�r2�����   ��3���]����������������������������������������������������������������������������������������������������������������������������������������U��   ]�������U����E�    �E�E��   �� M��M��   �� U�U��} ��   �E�8 ��   �M��U��E��8csm�uD�M��yu;�U��z �t�E��x!�t�M��y"�u�U��z u������   �E��M��QR�E�P�������E�����M􋐈   �����M����   ��u���M����   ��U�������E�� �����S���   �E�M����E��9�����    }�+��ǀ�       �   ��]���������������������������������������������������������������������������������������������U����E�E��   �� M��M��   �� U��U��E��8��G  �M�Q�s������} ��   �m�����   �:csm�u~�Z�����   �xum�I�����   �y �t(�5�����   �z!�t�!�����   �x"�u1������   �QR�#������tj�������   P�������������   �9csm�um�������   �zu\������   �x �t(������   �y!�t������   �z"�u �} t�v���   �E�E����U�
�\���M�����   �L���M�����   ��]��������������������������������������������������������������������������������������������������U����E��M�U��E��}�RCC�t(�}�MOC�t�}�csm�t�@���ǀ�       ����������    ~����   �E��M�����E��3��3���]����������������������������������������U��j�hp�h�Ld�    P���SVW���1E�3�P�E�d�    �e�E�x�   �M�Q���   �E��	�M�Q�U��E��E������   �E܋M܋���E܉�E�    �M�;M��   �}��~�U�E�;B}���1���M�Q�E�M��E�   �U�B�M�|� t%�U�E؉Bh  �MQ�U�B�M�T�R�5���E�    ��E�P��$����Ëe��E�    �M؉M��f����E������   �)������    ~�����   �EԋUԋ���MԉËU�;Uu��1���E�M�H�M�d�    Y_^[��]���������������������������������������������������������������������������������������������������U����E�     �H�����   �M��}� ��   �U��B�E��}� t%�M����t�E��H��U�E���E�M��R�U��B���E�M��Q��E���M����M��U���U�}� ~�E��M�U���t�M�   ���3���]������������������������������������������������U����q�����   u<�E�8csm�t1�M�9&  �t&�U�%���="�r�M�Q ��t
�   �  �E�H��ft4�U�z t�} uj��EP�MQ�UR��������   ��   ��   �E�x u$�M��������!���   �E�x ��   �M�9csm�uo�U�zrf�E�x"�vZ�M�Q�B�E��}� tH�M�Q� "������t1�U$R�E P�MQ�UR�EP�MQ�UR�EP�U��� �E��E��7��u.���)�M Q�UR�E$P�MQ�UR�EP�MQ�UR������ �   ��]���������������������������������������������������������������������������������������������������������U��Q�E�x t�M�Q�   k� �T
��u
�   �   �E���   t�U���t
�   �   �M�U�A;Bt$�M�Q��R�E�H��Q�a������t3��O�U���t
�M���t1�E���t
�U���t�M���t
�E���t	�E�   ��E�    �E���]�������������������������������������������������������������U�������E��E��Hl�M��U�;4�t�E��Hp# �u����E��U����   ��]����������������������������U���]�������U��Q�}�   s	�E�   ��E�    �E���]�������������U��Q�EP��-������u�M��_t	�E�    ��E�   �E���]����������������������������U��Q�EP��,������u�}_t	�E�    ��E�   �E���]����������������U��E��]������U����EP�M�������M��	-����t/�M���,����yt~�M���,��Ph  �UR��������E��h  �EP�M���,��P�������E��M��M��M������E���]����������������������������������U����EP�M��#����M��i,����t/�M��],����yt~�M��M,��Ph  �UR�6������E��h  �EP�M��%,��P��������E��M��M��M������E���]����������������������������������U����EP�M������}	u	�E�@   �X�M��+����t,�M��+����yt~�M��+��Pj@�UR�������E��j@�EP�M��|+��P�J������E��M��M��U��U�M��X����E��]���������������������������������������������������U����EP�M�������M��	+����t,�M���*����yt~�M���*��Pj �UR��������E��j �EP�M���*��P�������E��M��M��M������E���]����������������������������������������U��Q�EP�MQ�e�������u�}_t	�E�    ��E�   �E���]����������������������������U��Q�EP�MQ��������u�}_t	�E�    ��E�   �E���]����������������������������U����EP�M������M���)����t,�M��)����yt~�M��)��Pj�UR�������E��j�EP�M��)��P�Y������E��M��M��M��m����E���]����������������������������������������U����EP�M�������M��))����t/�M��)����yt~�M��)��Ph  �UR��������E��h  �EP�M���(��P�������E��M��M��M�������E���]����������������������������������U����EP�M��C����M��(����t,�M��}(����yt~�M��m(��Pj�UR�Y������E��j�EP�M��K(��P�������E��M��M��M��-����E���]����������������������������������������U����EP�M������M���'����t/�M���'����yt~�M���'��PhW  �UR�������E��hW  �EP�M��'��P�s������E��M��M��M������E���]����������������������������������U����EP�M������M��I'����t,�M��='����yt~�M��-'��Pj�UR�������E��j�EP�M��'��P��������E��M��M��M�������E���]����������������������������������������U����EP�M��c����M��&����t,�M��&����yt~�M��&��Pj�UR�y������E��j�EP�M��k&��P�9������E��M��M��M��M����E���]����������������������������������������U����EP�M�������M��	&����t,�M���%����yt~�M���%��Pj�UR��������E��j�EP�M���%��P�������E��M��M��M������E���]����������������������������������������U����EP�M��#����M��i%����t/�M��]%����yt~�M��M%��Ph�   �UR�6������E��h�   �EP�M��%%��P��������E��M��M��M������E���]����������������������������������U��=� uh  �EP�#������j �MQ������]����������������U��=� uh  �EP��"������j �MQ������]����������������U��Q�=� u'�}	u	�E�@   �j@�EP�"�����E��E���j �MQ��������]���������������������������U��=� uj �EP�9"������j �MQ�<�����]�������������������U��=� uj�EP��!������j �MQ������]�������������������U��=� uh  �EP�!������j �MQ������]����������������U��=� uj�EP�y!������j �MQ�W����]�������������������U��=� uhW  �EP�6!������j �MQ�X�����]����������������U��=� uj�EP�� ������j �MQ�/�����]�������������������U��=� uj�EP� ������j �MQ�"�����]�������������������U��=� uj�EP�y ������j �MQ������]�������������������U��=� uh�   �EP�6 ������j �MQ������]����������������U��j j j�EP�>����]����������U����E�    �} u3��l�EP�$��������E��MQ�UR�EPj�M�Q��������E��}� t5j jRh��hD�h`��UR�E�P�M�Q�H����P��������E��3���]������������������������������������������U����!���E��E��Hl�M��U�;4�t�E��Hp# �u����E��U��B��]�������������������������������U��������E��E��Hl�M��U�;4�t�E��Hp# �u�>���E��U��B��]�������������������������������U����a���E��E��Hl�M��U�;4�t�E��Hp# �u�����E��E��   ��]�����������������������������U�������E��E��Hl�M��U�;4�t�E��Hp# �u�~���E��U��Bt��]�������������������������������U��Q�} u
�d���E���E��Qt�U��E���]�����������U���@���3ŉE��E�    �E�    �E�    �E�    �E�    �E�E��E�    �   ��U��
�    �-  �E�x u5�M��Qh  �   ��E���   Qj �U�R��������t�  j^h��jj�������E�jbh��jjh�  ��������E�jdh��jjh�  ��������E�jfh��jjh�  �������E�jhh��jjh  �������Eԃ}� t�}� t�}� t�}� t�}� u��  �E��     �MԉM��E�    �	�U����U��}�   }�E�M���U���U��ۍE�P�M�QR�L ��u�  �}�v�  �E�E�j �M�QRh�   �E��   Ph�   �Mԃ�Qh   �   ��E���   Qj �;	����$��u�?  j �U�BPh�   �M؁��   Qh�   �Uԃ�Rh   �   ���M���   Rj ������$��u��  �}�~u�E�E��	�M���M�   k� �M����tQ�   �� �M����t>�   k� �U��
�E��	�M����M�   �� �E��9M��U�U�� ���j �E�HQ�U܁�   Rh   �E�Pjj �������u�E  �   k�3��M�f��   k��M�� �   k��M�� �   ���E�� �   ���U��
 �}�~�E�E��	�M���M�   k� �M����t[�   �� �M����tH�   k� �U��
�E��	�M����M�   �� �E��9M�� �  �E��M�f��A   ���h�   �U܁�   R�E�P������j�MЁ�   Q�U�R������j�E�   P�M�Q�o������U���    ��   �E���   �����J��   3�u#j h�Yj h�   h��j���������u�j�U���   -�   P�b�����j�M���   ��   R�H�����j�E���   ��   Q�.�����j�U���   P�������M��   �U�Ẻ��   �M܁�   �U���   �E��   �M���   �UЁ   �E���   �M؁��   �U���   �E�MȉHtj�U�R������3���   j�E�P������j�M�Q������j�U�R�v�����j�E�P�h�����j�M�Q�Z������   �   �   �U���    tE�E���   �����Ju2�E���    w&hD�h�Yj h�   h��j�_�������u̋Uǂ�       �Eǀ�       �Mǁ�   8��Uǂ�   ���Eǀ�   @��M�At   3��M�3��������]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���,�} ~,�EP�MQ�  ���E�U�;U}�E���E��M�M�E�    �E�    �E�    �}$ u�U��H�M$�}( t	�E�	   ��E�   j j �UR�EP�M�Q�U$R� �E��}� u3��<  �}� ~W3�uS�����3��u���rD�M���Q��������t#h��  �U��DP�������P�U�����E���E�    �M��M���E�    �U܉U�}� u3���  �E�P�M�Q�UR�EPj�M$Q� ��u
�  �z  j j �U�R�E�P�MQ�UR� ������E��}� u
�P  �K  �E%   tK�}  t@�M�;M ~
�.  �)  �U R�EP�M�Q�U�R�EP�MQ��������u
�   ��   ��   �U��U�}� ~W3�uS�����3��u��rD�M���Q���������t#h��  �U�DP������P�*
�����E���E�    �M؉M���E�    �UԉU��}� u�~�|�E�P�M�Q�U�R�E�P�MQ�UR���������u�V�T�}  u+j j j j �E�P�M�Qj �U$R� �E��}� u�'�%�#j j �E P�MQ�U�R�E�Pj �M$Q� �E��}� t�U�R�i������E�P�]������E���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�E��M�M��U��U�E����E��}� t�M����t�E����E��֋E+E�����]������������������������U��Q�E��;Ev	�E�   ��E�    �E���]�����������U��} t�E�M��U���U�E]������������������U����EP�M�������M(Q�U$R�E P�MQ�UR�EP�MQ�UR�M�����P�`�����$�E��M�������E���]����������������������������U��Q�} t[�E���E�M��U��}���  u�EP�
�����3�}���  t*3�u&h��h�Yj h  h��j�@�������u̋�]����������������������������������������U��j�h؄h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�    �E�    �} ��   j j%hH�h��h��j"jh����EPj j �M�Q�������P������� j&hL�jj�U�R��������E܃}� u3���  j j)hH�h��h��j"jj��EP�M�Q�U�Rj �v�����P������ ��tj�E�P������3��r  �M�Q�UR��������E�j�E�P�������}� u3��D  �"����E̋M̋Ql�UċE̋Hh�M��E�    j jEhH�h��h �j"j�U�Rj �E�Pj j �M�Q�������P������� ��t3���  jHhL�j�U���R�~������E؃}� u3��  �   �� E؉E�j jOhH�h��h��j"j�M�Qj��U�R�E�P�M�Qj �S�����P�x����� ��tj�U�R������3��S  �EĉE�j��������E�    �M���U�|
 t�E���M�| uC�U���E�| u�M���U�|
 t#hx�h�Yj jYhH�j�u�������u̋M���U�|
 t/�E���M�T�����Huj�M���U�D
P��������M̋Qp��uI� ���u?�M���U�|
 t/�E���M�T�����Huj�M���U�D
P�}������M؋U���M���U�E؉D
�M���U�EԉD
�E������   �j�������ËEԋM�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�   ��E�    �E��E܃}� u#hp�h�Yj j6h��j�"�������u̃}� u-�c���    j j6h��h��hp��������3��  �} t	�E�   ��E�    �U؉Uԃ}� u#h�h�Yj j7h��j調������u̃}� u-�����    j j7h��h��h��H�����3��  �M���t	�E�   ��E�    �EЉẼ}� u#h0�h�Yj j8h��j�.�������u̃}� u-�o���    j j8h��h��h0��������3��   ������E�}� u�4���    3��t�E�    �U���u*����    �E�    j��M�Qh���������E��9�U�R�EP�MQ�UR�������E��E������   ��E�P������ËEȋM�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������U��j@�EP�MQ�*�����]����������U����} t	�E�   ��E�    �E��E��}� u&h`�h�Yj h�   h��j�W�������u̃}� u0����    j h�   h��h��h`���������   �-h�   �UR�EP�������M��U�: t3���B��� ��]������������������������������������������������������������U����E�E��M��Q��   u�����    ����   �E��H���U��J�}u�E�P������E�E�E    �M�Q�������U��B%�   t�M��Q����E��P�-�M��Q��t"�E��H��t�U��B%   u
�M��A   �UR�EP�M�Q�`�����P����������u	�E�������E�    �E���]����������������������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h �h�Yj jch��j�	�������u̃}� u.�J���    j jch��h �h ������������   �} t�}t�}t	�E�    ��E�   �U܉U؃}� u#hȫh�Yj jdh��j脺������u̃}� u+�� ���    j jdh��h �hȫ�"���������H�MQ�������E�    �UR�EP�MQ��������E��E������   ��UR�?�����ËEԋM�d�    Y_^[��]�����������������������������������������������������������������������������������������������������U��j@�EP�MQ������]����������U����} t	�E�   ��E�    �E��E��}� u&h`�h�Yj h�   h��j�'�������u̃}� u0�h����    j h�   h��h(�h`���������   �-h�   �UR�EP��������M��U�: t3������� ��]������������������������������������������������������������U��j�h8�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�   ��E�    �E��E܃}� u#hp�h�Yj j6h��j��������u̃}� u-�C����    j j6h��h�hp�������3��  �} t	�E�   ��E�    �U؉Uԃ}� u#h�h�Yj j7h��j芷������u̃}� u-������    j j7h��h�h��(�����3��  �M���t	�E�   ��E�    �EЉẼ}� u#h0�h�Yj j8h��j��������u̃}� u-�O����    j j8h��h�h0�������3��   ������E�}� u�����    3��t�E�    �U���u*������    �E�    j��M�Qh��������E��9�U�R�EP�MQ�UR�n������E��E������   ��E�P�~�����ËEȋM�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������U����E�T=  �E�    �   k�����3���U�tj �E�P�U��E��}�zu�   �3���]���������������������U��Q�   k�����3���U�t�EP�U���]�������������������������U��Q�   k�����3���U�t�EP�U���]�������������������������U��Q�   k�����3���U�t�EP�MQ�UR�EP�U���MQ�U��R�E��P�MQ�` ��]�������������������������������U��Q�   k�����3���U�t�EP�MQ�UR�EP�MQ�UR�U���EP�MQ�UR�EP�� ��]�����������������������������U��Q�   k�����3���U�t�EP�MQ�UR�U��
jx�X 2���]���������������������U��Q�   ������3���M�t�UR�EP�MQ�U��3���]�����������������������������U��Q�   k�����3���U�t�EP�MQ�UR�U��3���]�����������������������������U��Q�   k� ����3���U�t	�EP�U���p ��]�����������������U��Q�   �� ����3���M�t	�UR�U��
�EP�| ��]�����������������������������U��Q�   ������3���M�t	�UR�U��
�EP�t ��]��������������U��Q�   k�����3���U�t�EP�MQ�U���UR�EP�x ��]���������������������U��Q�   k�����3���U�t�U���]�������������U��Q�   ������3���M�t�UR�EP�U���]���������������������U��Q�   k�����3���U�t�U��3���]�������������������������U��Q�   k�����3���U�t�EP�MQ�UR�EP�U��
jx�X 3���]�����������������U��Q�   k�����3���U�t�EP�MQ�U��
jx�X 3���]�������������������������U���H�E�P�� �M��t	�U�U���E�
   f�E���]�����������������U��Q�   k�����3���U�t�U���� 3ҋ�]�������������������U��Q�   ������3���M�t�UR�EP�MQ�U���UR�EP�\ �   ��]����������������������������U��Q�=� }
��������=� ~	�E�   ��E�    �E���]��������������������������U��Qh@��� �E�h`��E�P�� 3���   k� ����hl��E�P�� 3���   �� ����hx��U�R�� 3���   �ቁ��h���U�R�� 3���   k�����h���E�P�� 3���   ������h���U�R�� 3���   k�����h���E�P�� 3���   k�����h���E�P�� 3���   k�����h��E�P�� 3���   ������h ��U�R�� 3���   k�	����h8��E�P�� 3���   k�
����h`��E�P�� 3���   k�����h|��E�P�� 3���   k�����h���E�P�� 3���   k�����h���E�P�� 3���   k�����h���E�P�� 3���   k�����h���E�P�� 3���   ������h��U�R�� 3���   k�����h0��E�P�� 3���   k�����hX��E�P�� 3���   k�����hp��E�P�� 3���   k�����h���E�P�� 3���   k�����h���E�P�� 3���   k�����h���E�P�� 3���   k�����h���E�P�� 3���   k�����h���E�P�� 3���   k�����h���E�P�� 3���   k�����h��E�P�� 3���   k�����h0��E�P�� 3���   k�����h@��E�P�� 3���   k�����hX��E�P�� 3���   k�����hl��E�P�� 3���   k�����h���E�P�� 3���   ��������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�   ������3���M�t�UR�EP�MQ�UR�U��
jx�X 3���]�����������������U��Q�   k�����3���U�t	�EP�U��3���]���������������������U��Q�   k�	����3���U�t�EP�MQ�UR�EP�U���]�����������������������������U��Q�   k�����3���U�t�EP�MQ�UR�U���]�����������������U��EP�T ]������������������U��EP�d ]������������������U��EP�h P�l ]�����������U��j �T �EP�P ]����������U��Q�   k�
����3���U�t�EP�MQ�U���]���������������������U��Q���E��M��#M��U#Uʉ��E���]������������������������U��Q�E�    ����t
j
�D����������E��}� t
j�>���������t#j�o�����t�   �)jh  @j������j������]���������������������������������U���Ph��  h?  �������E��E%�  =�  ��   ���E�$�~������E��}� ~R�}�~�}�t�Dh��  �M�Q�j������E�j  �U�R�E�]��E؃��$���E�$j�������?  �E�P�E��`���$�E�]��EЃ��$���E�$jj�O�����$�  �E��������Dzh��  �M�Q��������E��  �U�R���E�$�������]�} }!�   �+E9E�}	�E�   ��	�M�M�M������+U9U�~	�E�����	�E�E�E��}� 
  ~M�M�Q���E��$���p��$�������$�E�]��Eȃ��$���E�$jj�t�����$�(  �}�   ~T�U���   R���E��$�w������]��E�P���E��$�E�]��E����$���E�$jj������$��   �}����}<�M�Q�E��x^���$�E�]��E����$���E�$jj�ң����$�   �}����}Q�U���   R���E��$�ս�����]��E�P���E��$�E�]��E����$���E�$jj�u�����$�,�M�Q���E��$芽�����]�h��  �U�R��������E���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�E��M�Q�UR�@�������]�������������������U��Q�E�E��M�Q�UR�EP讟������]���������������U��Q�E�E��M�Q�UR葟������]�������������������U��Q�E�E��M�Q�UR�EP�`�������]���������������U��Q�E�E��M�Qj �UR�EP�MQ�UR��������]���������������������U��Q�E�E��M�Q�UR�EP�MQ�UR�EP�T�������]�������������������U��Q�E�E��M�Q�UR�EP�MQ�v�������]�����������U��Q�E�E��M�Qj �UR�EP�MQ��������]�������������������������U��Q�E�E��M�Q�UR�EP�MQ�UR�h�������]�����������������������U��Q�E�E��M�Q�UR�EP�MQ�UR��������]�����������������������U���D�E�    3��E��EĉEȉẺEЉEԉE؍M��M��} t	�E�   ��E�    �U��U�}� u#h��h�Yj jih��j覠������u̃}� u.������    j jih��hD�h���D���������  �} t	�E�   ��E�    �M��M�}� u#hX�h�Yj jnh��j�-�������u̃}� u.�n����    j jnh��hD�hX������������   �E�E��M��A����U��BB   �E��M�H�U��E��M�Qj �UR�E�P��������E�} u�E��Q�M��Q���U�E��M�H�}� |"�U���  3Ɂ��   �M܋U�����M����U�Rj �������E܋E��]�����������������������������������������������������������������������������������������������������������������U��Q�E�E��M�Qj �UR�EP�MQ��������]������������������������̋T$�L$��   u@�:u2��t&:au)��t��:Au��t:au������uҋ�3���������Ë���   t���:u����t���   t�f���:u΄�t�:auń�t����������������������������������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^����������������������������U���������E��E��Hl�M��U�;4�t�E��Hp# �u�N����E�� ���]��������������������������������U��Q�����E��}� u	������E�����]������������U��V�C����M��UR����������0����0^]�����������U��Q�#����E��}� u	������E�����]������������U����} t	�E�   ��E�    �E��E��}� u&h��h�Yj h�   h��j�W�������u̃}� u%j h�   h��h �h����������   ��n����U� �3���]��������������������������������������U����} t	�E�   ��E�    �E��E��}� u&h��h�Yj h�   h��j觛������u̃}� u%j h�   h��h�h���M������   �������U� �3���]��������������������������������������U��Q�E�    �	�E����E��}�-s�M��U;͐�u�E��Ŕ��7�ԃ}r�}$w	�   �"� �}�   r�}�   w	�   ���   ��]�������������������������������U��Q�����E��}� u	�   ���ܟ���M�3���]����������������������U��Q������E��}� u	�   �������M�3���]����������������������U��j�hXd�    P�����3�P�E�d�    �EP�M��ģ���E�    �M�M�M�������P�E�L#Mu;�} t�M����������   �M�H#U�U���E�    �}� u	�E�    ��E�   �E�E��E������M�葳���E�M�d�    Y��]�������������������������������������������������U��jh  �EPj �������]�������U��jh  �EP�MQ�������]���������������������U��jh  �EPj ������]�������U��jh  �EP�MQ������]���������������������U��Q�}	u	�E�@   �jj@�EPj �N������E��E���]������������������U��Q�}	u	�E�@   �jj@�EP�MQ�������E��E���]����������������U��jh  �EPj �������]�������U��jh  �EP�MQ������]���������������������U��jj �EPj ������]����������U��jj �EP�MQ�l�����]��������U��j �EP�m�����]��������������U����EP�M��#����M��i����x t8�M��[����H�y�  u$jj �UR�EP��������E��M��,����E���E�    �M������E���]�����������������������������������U��jj �EPj ������]����������U��jj �EP�MQ�|�����]��������U��jj �EPj �^�����]����������U��jj �EP�MQ�<�����]��������U��jj �EPj ������]����������U��jj �EP�MQ�������]��������U��jhW  �EPj �������]�������U��jhW  �EP�MQ������]���������������������U��jj�EPj ������]����������U��jj�EP�MQ�l�����]��������U��jj �EPj �N�����]����������U��jj �EP�MQ�,�����]��������U����E�E��M���U��E����E��}� t��E�+E������]����������������������������U��j �q�����]������������������U���(V�E�    �EP�M�苞���M����������   �U��E�    �	�E����E��}�s3�M��U��P踾�������M��U�D�P裾����E�L0�M��jChD�j�U��R�q������E��}� ��   �E��E��E�    �	�M����M��}���   �U��:�E����E�j jJhx�h��h���M��U��P�M���U�+U�+�Q�E�P�d�����P袞�����M�Q�������E��E��U��:�E����E�j jMhx�h��hx��M��U�D�P�M���U�+U�+�Q�E�P������P�?������M�Q葽����E��E��#����U�� �E����E��M��M�M��I����E�^��]�������������������������������������������������������������������������������������������������������������������U��j ������]������������������U���(V�E�    �EP�M��K����M���������   �U��E�    �	�E����E��}�s4�M��U�D�8P�w��������M��U�D�hP�b�����E�L0�M��jjhD�j�U��R�0������E��}� ��   �E��E��E�    �	�M����M��}���   �U��:�E����E�j jqhx�h��h��M��U�D�8P�M���U�+U�+�Q�E�P�"�����P�`������M�Q費����E��E��U��:�E����E�j jthx�h��h���M��U�D�hP�M���U�+U�+�Q�E�P������P��������M�Q�O�����E��E��"����U�� �E����E��M��M�M������E�^��]�����������������������������������������������������������������������������������������������������������������U��j �v�����]������������������U��j �EP�MQ�UR�EP�MQ词����]��������������U���T�E�    �E�    �E�    �EP�M��Ι���} t	�E�   ��E�    �M�M�}� u&h��h�Yj h�   hx�j�Ə������u̃}� u@�����    j h�   hx�h(�h���a������E�    �M�蒩���E��  �} t	�E�   ��E�    �E�E��}� u&hD�h�Yj h�   hx�j�8�������u̃}� u@�y����    j h�   hx�h(�hD���������E�    �M������E��  �U� �} t	�E�   ��E�    �E܉E؃}� u&hl�h�Yj h�   hx�j褎������u̃}� u@������    j h�   hx�h(�hl��?������E�    �M��p����E���  �} t	�E�   ��E�    �UԉUЃ}� u&h��h�Yj h   hx�j��������u̃}� u@�W����    j h   hx�h(�h���������E�    �M������E��^  j j j��MQj �M��������BP� �E��}� u�� P�f�������   h
  hD�j�M���Q蕉�����E��}� u��   �U�R�E�Pj��MQj �M��a�����BP� ��u�� P�������   h  hD�j�M��Q�1������E��}� u�k�UR�EP�MQ�U�R�EP�M�Q�d������E�}� tBj j �UR�EPj��M�Qj �M��������BP� ��u�� P�t������E�    j�M�Q�,�����j�U�R�������E�E��M������E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP�MQ迈����]��������������U��j j �EP�MQ�UR�EP葈����]����������������U���   V�E�E��M����M��}�v��  �U�����$����M�y |�U�zǅl���   �
ǅl���    ��l����E�}� u&h��h�Yj h�  h �j胊������u̃}� u0������    j h�  h �h,�h��������3��X  �UR�EP�M�Q�E����   Q�  ���-  �U�z |�E�x	�E�   ��E�    �M��M܃}� u&h��h�Yj h�  h �j�Ӊ������u̃}� u0�����    j h�  h �h,�h���n�����3��  �EP�MQ�U�B�M����   R�j  ���}  �E�x |�M�yǅ\���   �
ǅ\���    ��\����Uԃ}� u&hP�h�Yj h�  h �j��������u̃}� u0�[����    j h�  h �h,�hP�������3���  �MQ�UR�E�H�U����   P�  ����  �M�y |�U�z	�E�   ��E�    �E��Ẽ}� u&hP�h�Yj h�  h �j�j�������u̃}� u0�����    j h�  h �h,�hP�������3��?  �UR�EP�M�Q�E���  Q�  ���  �}  ��   �UR�EP�MQ�URj�EP�4  ����u3���  �M�9 u3���  �U��    f��U����M��U����M��UR�EP�MQ�URj�EP��  ����u3��  �   �MQ�UR�EP�MQj �UR�  ����u3��Y  �E�8 u3��J  �M��    f��M����E��M����E��MQ�UR�EP�MQj�UR�H  ����u3���  ��  �E�x|�M�yǅt���   �
ǅt���    ��t����Uă}� u&h��h�Yj h(  h �j荆������u̃}� u0������    j h(  h �h,�h���(�����3��b  �M Q�UR�EPj�M�QR�h  ���;  �E�x |�M�y	�E�   ��E�    �U��U��}� u&hh�h�Yj h1  h �j��������u̃}� u0�"����    j h1  h �h,�hh��|�����3��
  �M Q�UR�EPj�M�QR�  ���
  �E�x |�M�yǅd���   �
ǅd���    ��d����U��}� u&hh�h�Yj h9  h �j�,�������u̃}� u0�m����    j h9  h �h,�hh��������3��
  �M�A��   ���U��}� u�E�   �U R�EP�MQj�U�R��  ���	  �E�x |�M�ym  	�E�   ��E�    �U��U��}� u&h��h�Yj hD  h �j�b�������u̃}� u0�����    j hD  h �h,�h���������3��7	  �M Q�UR�EPj�M�Q��R�:  ���	  �E�x |�M�y	�E�   ��E�    �U�U��}� u&hP�h�Yj hM  h �j賃������u̃}� u0������    j hM  h �h,�hP��N�����3��  �M Q�UR�EPj�M�Q��R�  ���^  �E�x |�M�y;ǅ|���   �
ǅ|���    ��|����U�}� u&h� h�Yj hV  h �j���������u̃}� u0�<����    j hV  h �h,�h� ������3���  �M Q�UR�EPj�M�QR��  ���  �E�x |�M�y	�E�   ��E�    �U��U؃}� u&hh�h�Yj h^  h �j�O�������u̃}� u0�����    j h^  h �h,�hh��������3��$  �M�y%�UR�EP�   k� �E��L  Q��  ���#�UR�EP�   �� �U��
L  P�  ����  �M�9 |�U�:;	�E�   ��E�    �EЉEȃ}� u&hh�Yj hi  h �j�q�������u̃}� u0�����    j hi  h �h,�h������3��F  �U R�EP�MQj�U�P�M  ���   �M�y |�U�z	�E�   ��E�    �E��E��}� u&h��h�Yj hp  h �j�ƀ������u̃}� u0�����    j hp  h �h,�h���a�����3��  �U�B�E��Y  �T  �M�y |�U�z	�E�   ��E�    �E��E��}� u&h��h�Yj hw  h �j�)�������u̃}� u0�j����    j hw  h �h,�h���ľ����3���  �U R�EP�MQj�U�BP�
  ����  �M�y |�U�z	�E�   ��E�    �E��E��}� u&h��h�Yj h~  h �j�}������u̃}� u0�����    j h~  h �h,�h��������3��R  �U�z u	�E�   ��E�H���M�U�z |�E�xm  	�E�   ��E�    �M��M��}� u&h��h�Yj h�  h �j��~������u̃}� u0�����    j h�  h �h,�h���m�����3��  �E�H;M�}	�E�    �-�U�B��   ���E��U�B��   ��;U�|	�U����U��E P�MQ�URj�E�P�o  ���B  �}  t+�MQ�UR�EP�MQj�UR�f
  ����u3��  �)�EP�MQ�UR�EPj �MQ�;
  ����u3���  ��  �UR�EP�MQ�URj�EP�
  ����u3��  �  �M�y |	�E�   ��E�    �U���x�����x��� u&h�h�Yj h�  h �j�^}������u̃�x��� u0�����    j h�  h �h,�h��������3��0  �M�A��d   ���U��U R�EP�MQj�U�R�(  ����  �E�x����|�M�y�  ǅp���   �
ǅp���    ��p�����h�����h��� u&h�h�Yj h�  h �j�|������u̃�h��� u0������    j h�  h �h,�h��$�����3��^  �M�A��d   ����k�d�U�B��d   ��ʉM��E P�MQ�URj�E�P�@  ���  ������E�    �M�y  tǅ`���   �
ǅ`���    j h�  h �h,�hpj"j�URj��,�����`�����R�E�Q�U�P�M�Q�v�����P�y���� ��X�����X���Pu�U�    ��E����M�+ЋE��M��E��LB��U�
�Y�E��%   f��E����U�
�E����U�
�0�.3�u&hhh�Yj h�  h �j��z������u�3���   ^��]ÍI k�B�n�ל`��=�ң{�ĥ�������������ܠ����Y��m�  	
���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�    �} t�EP�MQ�UR�   ���   �E�M;sn�U���U�	�E���E�M��t3�E��
   ����0�E��Ef�A�E��
   ���E�U����U�뼋E��U��Q�M��U�+E��M��	�U�    ��]��������������������������������������������������U����E��M��U�:vF�E��
   ����0�E�f��M����M��U����M��E��
   ���E�} ~�U�:w��E��M�U�E���M����M��U�f�f�E��M��U�f�f��M����M��U�f�E�f��M���M�U�;U�rƋ�]����������������������������������������������U��E�8 t=�M���t3�E��Uf�f��M����E��M���M�U����M��]�����������������������U���h���3ŉE��E�E��}� t�}�t��M��T  �U���E��X  �M���U��\  �E�M���   ��  �E�   �}t�E�    �U�Bl  f�E�M�Q��f�U�Ef�Hf�M�Uf�Bf�E�Mf�Qf�U��Ef�f�M�3�f�U��}� t%j j �E�P�M�Qj �U��`  P�s������E��#j j �M�Q�U�Rj �E��`  Q�>������E؃}� �  �U���R��~������t#h��  �E؍L Q跜����P�7������E���E�    �U��Ũ}� ��   �}� t)�E�P�M�Q�U�R�E�Pj �M��`  R�˄�����E��'�E�P�M�Q�U�R�E�Pj �M��`  R蒲�����E؋ẺE܋M؃��M؃}� ~;�U�: v3�E��U�f�f��M����E��M܃��M܋U����M�붋U�R�a������   �  �E������  �U�: ��  3�f�E��E�    �E�    �M�M��	�U����U��E���M��U���E��M܃��M܋U�;U�u�ҋE܃��E܋M���UċEă�'�Eă}�R�
  �M���D��$���E��E��M����M��}�w0�U��$����E�   �m   f�E���b   f�M��	�B   f�U��  �E��EȋMȃ��Mȃ}�w0�U��$����E�   �d   f�E���a   f�M��	�A   f�U��e  �E��E��}�t�}�t��y   f�M��	�Y   f�U��8  �E��E��}�t�}�t	��E�   �I   f�M��  �U��U��}�t�}�t	��E�   �H   f�E���  �M��M��}�t�}�t	��E�   �M   f�U��  �E��E��}�t�}�t	��E�   �S   f�M��  h��U�R輅������u�E��
�E��h��M�Q蜅������u	�U���Uܸp   f�E��H  �M�y�   k� �M��L  �U���   �� �M��L  �Uԃ}�u;�E�8 v3�M��E�f�f�
�U����M��Uԃ��UԋE����U�
�E�E����t;�U�: v3�E��U�f�f��M����E��Mԃ��MԋU����M�뻋U܉U�������E���ti�M��U�J�E�M����tQ�E�8 tI�M����'u�E���E��3�M��E�f�f�
�U����M��U���U�E����U�
���E��M�A�U��m����E��t5�M�Q�UR�EP�MQ�UR�E�P�MQ���������u3��C�U܉U��1�E��U�f�f��M����E��M���M�U����M�������   �M�3��G�����]Ë���������X���ӵH�+��� 







































































	�����ȴӴ ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �Z�����]������������������U���(V�E�    �EP�M��t���M���������   �U��E�    �	�E����E��}�s:�M��U싄��   P�\��������M��U싄��   P�D�����E�L0�M��jHh��j�U�DP�f�����E��}� �  �M��M��E�    �	�U����U��}���   �:   �M�f��U����U�j jOh �hd�h���E��M싔��   R�E���M�+M���+�P�U�R������P�t�����E�P艓�����M��A�U��:   �M�f��U����U�j jRh �hd�h��E��M싔��   R�E���M�+M���+�P�U�R袰����P�?t�����E�P�������M��A�U�����3��M�f��U����U��E��E�M��D����E�^��]������������������������������������������������������������������������������������������������������������������������������U��j �p����]������������������U���(V�E�    �EP�M��;r���M�聵������   �U��E�    �	�E����E��}�s:�M��U싄��   P���������M��U싄�  P�ԑ����E�L0�M��joh��j�U�DP�d�����E��}� �  �M��M��E�    �	�U����U��}���   �:   �M�f��U����U�j jvh �h��h���E��M싔��   R�E���M�+M���+�P�U�R袮����P�?r�����E�P�������M��A�U��:   �M�f��U����U�j jyh �h��h8��E��M싔�  R�E���M�+M���+�P�U�R�2�����P��q�����E�P詐�����M��A�U�����3��M�f��U����U��E��E�M��Ԁ���E�^��]������������������������������������������������������������������������������������������������������������������������������U��j �6l����]������������������U���T�EP�M���o���M���������   �U��E�    �E�d  �E�    �E�    �	�E����E��}���  �}�uWh�   h��j�M�Q��a�����E��}� u�E�    �M�����E��  �U�Rj �E�P莌�����M��M��E�d  �E�    �	�U���U�}���   �E�3ҹ   ���t�U����U���}�uQ�E�E��M�U���j h�   h �h��h���E�M��R�E�+E�P�M�U���P�r�����P�o�����M�U��P��������M��T�U��Z����E�    �	�E���E�}���   �E�3ҹ   ���t�U����U���}�uT�E�E��M�U��D�j h�   h �h��h���E�M�T�R�E�+E�P�M�U��D�P�������P��n�����M�U�D�P�I������M��T�U��V����E�    �	�E����E��}���   �E�3ҹ   ���t�U����U���}�uT�E�E��M��U��D�8j h�   h �h��hp��E��M�T�8R�E�+E�P�M��U��D�8P������P�Kn�����M��U�D�8P薍�����M��T�U��V����E�    �	�E܃��E܃}���   �E�3ҹ   ���t�U����U���}�uT�E�E��M܋U��D�hj h�   h �h��hP��E܋M�T�hR�E�+E�P�M܋U��D�hP�Z�����P�m�����M܋U�D�hP�������M��T�U��V����E�    �	�E؃��E؃}���   �E�3ҹ   ���t�U����U���}�u]�E�E��M؋U�����   j h�   h �h��h��E؋M􋔁�   R�E�+E�P�M؋U�����   P螩����P��l�����M؋U􋄊�   P�$������M��T�U��J����E�3ҹ   ���t�U����U���}�uQ�E�E��M����   j h�   h �h��h���U􋂠   P�M�+M�Q�U����   P������P�El�����M􋑠   R葋�����M��T�U��E�3ҹ   ���t�U����U���}�uQ�E�E��M����   j h�   h �h��h���U􋂤   P�M�+M�Q�U����   P�y�����P�k�����M􋑤   R�������M��T�U��E�3ҹ   ���t�U����U���}�uQ�E�E��M����   j h�   h �h��hx��U􋂨   P�M�+M�Q�U����   P������P�)k�����M􋑨   R�u������M��T�U��}�u�E��M􋑬   ���   �E�ǀ�       �E�    �	�Mԃ��Mԃ}���   �E�3ҹ   ���t�U����U���}�ud�E���M��A�EԋM�����   j h�   h �h��h@��UԋE􋌐�   Q�U�+U���R�EԋM�����   R誦����P�Gj�����EԋM􋔁�   R�������M��TA�U��C����E�    �	�EЃ��EЃ}���   �E�3ҹ   ���t�U����U���}�ud�E���M��A�EЋM�����   j h�   h �h��h0��UЋE􋌐�   Q�U�+U���R�EЋM�����   R������P�i�����EЋM􋔁�   R�Q������M��TA�U��C����E�    �	�Ẽ��Ẽ}���   �E�3ҹ   ���t�U����U���}�ud�E���M��A�E̋M�����   j h�   h �h��h��ŰE􋌐�   Q�U�+U���R�E̋M�����   R������P�h�����E̋M􋔁�   R苇�����M��TA�U��C����E�    �	�Eȃ��Eȃ}���   �E�3ҹ   ���t�U����U���}�ud�E���M��A�EȋM����  j h�   h �h��h ��UȋE􋌐  Q�U�+U���R�EȋM����  R�X�����P��g�����EȋM􋔁  R�ņ�����M��TA�U��C����E�    �	�Eă��Eă}���   �E�3ҹ   ���t�U����U���}�ud�E���M��A�EċM����L  j h�   h �h��h���UċE􋌐L  Q�U�+U���R�EċM����L  R蒣����P�/g�����EċM􋔁L  R��������M��TA�U��C����E�3ҹ   ���t�U����U���}�uX�E���M��A�E���T  j h�   h �h��h���M�T  R�E�+E���P�M���T  R�������P�f�����E�T  Q�e������U��DB�E��E�3ҹ   ���t�U����U���}�uX�E���M��A�E���X  j h�   h �h��h���M�X  R�E�+E���P�M���X  R�_�����P��e�����E�X  Q�Є�����U��DB�E��E�3ҹ   ���t�U����U���}�uX�E���M��A�E���\  j h�   h �h��hx��M�\  R�E�+E���P�M���\  R�ʡ����P�ge�����E�\  Q�;������U��DB�E��E�3ҹ   ���t�U����U���}�uX�E���M��A�E���`  j h�   h �h��hX��M�`  R�E�+E���P�M���`  R�5�����P��d�����E�`  Q覃�����U��DB�E������M��M��M���s���E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�EP�MQ�r����]��������������U���l�E�    �E�E��MQ�M��&`���} t	�E�   ��E�    �U�U��}� u&h��h�Yj h  h �j�V������u̃}� u@�_����    j h  h �hH�h��蹔�����E�    �M���o���E��  �} t	�E�   ��E�    �M�M�}� u&hD�h�Yj h  h �j�U������u̃}� u@�ћ���    j h  h �hH�hD��+������E�    �M��\o���E��   3��Mf��} t	�E�   ��E�    �U�U��}� u&hl�h�Yj h  h �j��T������u̃}� u@�;����    j h  h �hH�hl�蕓�����E�    �M���n���E��j  �} u�M�贡������   �U���E�E܋M܉M��U�U��}� �N  �E��M؃}� t�}�%t
�  �/  �} t	�E�   ��E�    �UԉUЃ}� u&hd�h�Yj h7  h �j�T������u̃}� u@�W����    j h7  h �hH�hd�豒�����E�    �M���m���E��  �M���M�E�    �U���#u�E�   �M���M�U�R�E�P�M�Q�UR�EP�M�R�M�萠��P�g�������u�}� v�E�   �7�E���E�'�M�Uf�f��M���M�U���U�E����E������}� u,�}� v&3ɋUf�
�E+E��E��M��m���E��   �   3ɋU�f�
�}� u�}� w�0���� "   �v�E�    �}� u&h��h�Yj hw  h �j�R������u̃}� u=�����    j hw  h �hH�h���D������E�    �M��ul���E���E�    �M��al���E���M��Tl����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP�MQ�l����]��������������U��j j �EP�MQ�UR�EP�`l����]����������������U��E�� ]������U���<�EP�M��sZ���}   ��   �M�謝����t,�M�蠝����yt~�M�萝��Pj�UR�|d�����E��j�EP�M��n���P�<L�����E��}� t,�M��T�������   �E��M�M��6j���E��  ��U�U��M��j���E��  �M������ �xt~q�M�����P�M�����   Q��������tO�U�����   �   k� �T��   �� �E�D��   ��M�}�s��h����U��D� �E�   �=�ҕ��� *   �   k� �U�T��E�   �}�s��)����E��D� �E�   j�M��R�����QRj�E�P�M�Q�U�Rh   �M��1���� �   �ዔ�   R�M�����P������$�E�}� u�E�E܍M���h���E��\�}�u�   k� �D��E؍M���h���E��9�/�   �� �T��   k� �D���ЉUԍM��h���E���M��h����]�������������������������������������������������������������������������������������������������������������������������������������������������U��Q�=� u$�}A|�}Z�E�� �E���M�M��E���j �UR�v������]�����������������������������̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[����������������������������������������������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ����������������������������������������U����E�E��M�M��U���M��+�P�  ����]��������������������U��� �E�E��M�M�U�E��
;��   �U�U��E�E�M�Q�U�R�������E��}� t�E��E��s�M���Q�U��R�^������E��}� t�E��E��F�M���Q�U��R�7������E��}� t�E��E���M���Q�U��R�������E��E��E�M�M�E��3���]����������������������������������������������������U��Q�} t�} ~	�E�   ��E������E��E�E��]��������������������U����E�E�M�M�U���M��;�tK�E�E��M�M�U�R�E�P�E������E��}� t�M��M���U���R�E��P�������E��E��3���]������������������������������U���(�E�E��M�M�U�U��}��g  �E��$�$��M�Q�U�R�������E��}� t�E��E��s�M���Q�U��R�������E��}� t�E��E��F�M���Q�U��R�i������E��}� t�E��E���M���Q�U��R�B������E�E�E�M�M�E���   �U�R�E�P�������E��}� t�M��M��F�U���R�E��P��������E��}� t�M��M���U���R�E��P��������E��M��M܋E��i�U�R�E�P�������E��}� t�M��M���U���R�E��P�������E؋E��*�M�Q�U�R�p������3���EP�M�Q�U�R�   ����]ÍI �����H���������������������������������������������������������������������������������������������������������������������������U����} �R  �EP�MQ��������E��}� t�E��O  �U��R�E��P�������E��}� t�E��(  �M��Q�U��R�������E��}� t�E��  �E��P�M��Q�n������E��}� t�E���  �U��R�E��P�G������E��}� t�E��  �M��Q�U��R� ������E��}� t�E��  �E��P�M��Q��������E��}� t�E��e  �U��R�E��P��������E��}� t�E��>  �M�� �M�U�� �U�E�� �E�����MM�M�UU�U�E�E��}���  �M��$�4��U��R�E��P�_������E��}� t�E���  �M��Q�U��R�8������E��}� t�E��  �E��P�M��Q�������E��}� t�E��}  �U��R�E��P��������E��}� t�E��V  �M��Q�U��R��������E��}� t�E��/  �E��P�M��Q�������E��}� t�E��  �U��R�E��P�u������E��}� t�E���  3���  �M��Q�U��R�G������E��}� t�E��  �E��P�M��Q� ������E��}� t�E��  �U��R�E��P��������E��}� t�E��e  �M��Q�U��R��������E��}� t�E��>  �E��P�M��Q�������E��}� t�E��  �U��	R�E��	P�������E��}� t�E���  �M��Q�U��R�]������E��}� t�E���  �E��P�M��Q��������  �U��R�E��P�������E��}� t�E��  �M��Q�U��R��������E��}� t�E��`  �E��P�M��Q��������E��}� t�E��9  �U��R�E��P�������E��}� t�E��  �M��Q�U��R�������E��}� t�E���  �E��
P�M��
Q�X������E��}� t�E���  �U��R�E��P�1������E��}� t�E��  �M��Q�U��R�J������  �E��P�M��Q��������E��}� t�E��[  �U��R�E��P��������E��}� t�E��4  �M��Q�U��R�������E��}� t�E��  �E��P�M��Q�z������E��}� t�E���   �U��R�E��P�S������E��}� t�E��   �M��Q�U��R�,������E��}� t�E��   �E��P�M��Q�������E��}� t�E��t�U��R�E��P�������E��}� t�M��M��F�U��R�E��P�z������E��}� t�M��M���U��R�E��P�S������E�M�M��E��3���]�O�g�����(�@�l�����E�q������J�������#���������e�}�����>�V���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���@���3ŉE��} ~�EP�MQ��  ���E��}�}3���  �}  ~�U R�EP��  ���E ��} �}3��  �E�    �}$ u�M��B�E$�} t
�}  ��  �M;M u
�   �o  �} ~
�   �_  �}~
�   �O  �U�R�E$P�L ��u3��6  �} u�} t2�}u�}  t&h�h�Yj h�   hpj�>������u̃} ��   �}�s
�   ��  �U�U��	�E���E�   k� �E����tQ�   �� �E����t>�U��   k� �M��;�|#�E��   �� �E��;�
�   �k  듸   �_  �}  ��   �}�s
�   �E  �E�E��	�M���M�   k� �M����tQ�   �� �M����t>�E��   k� �U��;�|#�M��   �� �M��;�
�   ��  듸   ��  j j �MQ�URj	�E$P� �E��}� u3��  �}� ~W3�uS�����3��u���rD�U���R��H������t#h��  �E��L Q�f����P�(~�����E���E�    �UЉU���E�    �E��E؃}� u3��'  �M�Q�U�R�EP�MQj�U$R� ��u
��   ��   j j �E P�MQj	�U$R� �E܃}� u
��   ��   �}� ~W3�uS�����3��u܃�rD�M���Q�H������t#h��  �U܍DP��e����P�\}�����E���E�    �MĉM���E�    �ỦUԃ}� u�Q�O�E�P�M�Q�U R�EPj�M$Q� ��t#�U�R�E�P�M�Q�U�R�EP�MQ��q�����EȋU�R��R�����E�P��R�����EȋM�3���Y����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�E��M�M��U��U�E����E��}� t�M����t�E����E��֋E+E�����]������������������������U����EP�M��CC���M$Q�U R�EP�MQ�UR�EP�MQ�M��m���P�D����� �E��M��US���E���]��������������������������������U����E�    �E��   �E�;E�A�E�E��+����E��M��U+�x�U�u�E���}� }�E����E��	�M����M�뷃����]�����������������������������U����E�X�E�    �E��   �E�;E�W�E�E��+����E�jU�M��U���P�MQ�4<�����E�}� u�U��E��D���}� }�M����M��	�U����U�롃����]������������������������������������������������U��Q�   k�����3���U�t#j j j �EP�MQ�UR�EP�MQ�UR�U��'�EP�MQ�UR�EP�MQ�UR�F����P�� ��]��������������������������������������U����} t�}   t	�}   u3��   �} u�} �} }3��   �EP�|R�����E��}� }3��i�M���|�U�jU�E�P�s�����E�} ~?�M�;M|3��9j h�   h -hd-h�-�U�R�EP�MQ��}����P�wA�����E����]�������������������������������������������������������������U��Q�} u3��,�EP�x�����E��}� |	�}��   r3��
�M���x��]�������������������U��j j �EP�\�]� �����������U����E�    �   k�����3���U�tj �EP�MQ�UR�U��%�E�\�jh���� �E��\�    �E���]�������������������������������U��Q�   k�����3���U�tj �EP�MQ�UR�EP�MQ�UR�U��'�EP�MQ�UR�EP�MQ�UR�C����P�� ��]��������������������������U��Q�   k�����3���U�t�EP�MQ�UR�EP�U���MQ�UR�EP�MQ�#C����P�� ��]����������������������������U��Q�   k�����3���U�t�EP�MQ�UR�EP�MQ�UR�U��'�EP�MQ�UR�EP�MQ�UR�B����P�� ��]����������������������������U��Q�   k�����3���U�t�EP�MQ�U���UR�EP�� P�VZ������]����������������������������U��Q�   k�����3���U�t	�EP�U��j�MQ��A����P�� ��]������������������U��Q�   k�����3���U�t#j j j �EP�MQ�UR�EP�MQ�UR�U��'�EP�MQ�UR�EP�MQ�UR�mA����P�� ��]��������������������������������������U����E�    �} ��   �E���A|�U���Z�M��� �U��	�E��M�f�U�f�U��E���A|�U���Z�M��� �U��	�E��M�f�U�f�U��E���E�M���M�U���Ut�E���t�M��U�;��a����E��M�+��E�E��]�������������������������������������������������������U����} ~�EP�MQ�un�����E�} ~�UR�EP�\n�����E�} t�} u4�M+Mu	�E�   ��U+Uy	�E�   ��E�   �E��E��E�� �MQ�UR�EP�MQ�UR�EP��g������]�����������������������������������������������������U��} ~�EP�MQ�m�����E�UR�EP�MQ�UR�EP�MQ�+����]�������������������U��j�h��h�Ld�    P��$SVW���1E�3�P�E�d�    �e��E� �E�  �E�EЍE�E��E�    �E�Pjj h�m@�8 ��E� 3Ɂ8�m@����Ëe��E������E�M�d�    Y_^[��]����������������������������������������U��j�h��h�Ld�    P��$SVW���1E�3�P�E�d�    �e��E� �E�  �E�EЋE�EԋE�E؍E�E܋E�E��E�    �E�Pjj h�m@�8 ��E� 3Ɂ8�m@����Ëe��E������E�M�d�    Y_^[��]������������������������������������������������������U���H  ���3ŉE��EW�=`��������E����������2  S�� Vh   j h`3�Ӌ���u"�� ��W��   VVh`3�Ӌ�����   h|3V�� �ȉ`�����   ����������   ����   �C�s h�3�u��$h�3Ph 4Vh,4h@4������h�4P�ыC��$PV�E�P�E�P�  ��8�E�h�4Ph�4�E�P������h�4P�  ��������P�`�������PjW�������  ��(^[_�M�3��~L����]�h�3jW��������  ��^[�M�3�_�WL����]�����������������������������������������������������������������������������������������������������������U��E��w#��P��� .���t.RPQ�u�7  ��]Ë4.�   RP�   Q�u�  ��]�����������������������������������U���  ���3ŉE��E�������X�������S�]�����   �; ��   S�  ��-��=   ��   3����$    ���P.�@��������u�VW��C��u�������+�O�GG��u��˺l.���˃���B��u�������+�O�GG��u��ʍ��������ʃ��_^��03Pj�������������  ���M�3�[�}J����]�����������������������������������������������������������������U��Q�U�MSVW�}3�+׉U�E�M���r�   ;�s%�:��Phd�Q�`��M����UF���G�ǋE_� �E�p� ^[��]�����������������������������������������U��U�@��u�+�H]�������������U���<  ���3ŉE��ES�]V�uWV������������ǅ����    �@M��������uV�D����������j j j�S� j h��  ��=   s#P������Pj�������j h��  �Ӎ�������u�2h  �~�������t$������SV�4�8.P�"��������  2��������� u����   ��t�  ����   h  ������P������Ph  ������P�F�P��h������t*S������������h�2P������������P�u���   � ������j j h
  Pj���������2Pj h��  �Ӆ�t������j j h
  ��������2Pj�������Pj h��  �Ӆ�t������������������h3V������W�u����������u̋M�_^3�[�G����]����������������������������������������������������������������������������������������������������������������������������������U���  ���3ŉE��\�������S�]�����   ����   S�7�����:��=   w3����    ���.�@��������u�VW��C��u�������+�O�GG��u��˺�.���˃���B��u�������+�O�GG��u��ʍ��������ʃ��_^���4P�Ej������P�������M�3�[�/F����]������������������������������������������������������������������̡d�����������̡h������������U��E��w	��5]�3�]��������̸   �����������U��d��M�d��h�    ]��������������������U��h��M�h��d�    ]��������������������U��U��w��P��M��P�]Ã��]��������������U���%]�������U�츌%]�������u�U��� PRSVWh�5h�Qj7h�6j�U&������u�_^[ZX��]�������������������������U��j��a������tj��a������u#�=p�uh�   �O����h�   �O����]����������������������������U��Q�E�    �	�E����E��}�s�M��U;�(7u�E���,7���3���]������������������U���   ���3ŉE��EP��.���������������� �  ǅ����    �}�   t\�}�   tS�}tM������Qh�Yj j j j�$���������������� t������t��ǅ����   �
ǅ����   ������ �  j�`������tj�`��������   �=p���   j��� ������������ ��   ���������   ǅ ���    ��� ������� ����� ����  s4�� ����� ����������J������� ����������P��u�뱺   i��  �������������  s��nb��������Ƅ��� j ������R�����P�M����P�����Q������R�� ��  �}�   ��  �   k���x�������������x����  +����������������j h  h�Bh Ch Ch�Ch  hx��j����P�-�����   i�  3ɋ����f�h  �����Pj �( ��u:j h  h�Bh Ch0Dh$�������Q�����R�i����P�G-����������P�L��������<vk�����Q�L�����������DB�������j h#  h�Bh Ch�Djh|�������+������������+�R������P�8����P��,����j h&  h�Bh ChXEh��h  hx���i����P�,����j h'  h�Bh Ch�E������Qh  hx��i����P�W,����h  h �hx��A�����M�3��.@����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE��}��  �E��h�����|�����x���ǅd���    ǅl����   ��l���R��x���P�MQ�UR�EP��i������p�����p��� ��   �� ��zt�/  j j �MQ�UR�EP�i������l�����l��� u�  j^h�Fjj��l���Q�8������x�����x��� u��   ǅd���   ��l���R��x���P�MQ�UR�EP�#i������p�����p��� u�   jih�Fjj��p���Q�7������h������h����8 u�fj jlh�Fh4Gh`G��p�����Q��x���R��p���P��h����R��j����P�)������d��� tj��x���P�]-����3��6  ��d��� tj��x���Q�<-��������  �  �}��   �U��t�����t����     j j �MQ�UR�l������`�����`��� u�\h�   h�Fjj��`���P�6������t������t����: u�*��`���P��t����R�EP�MQ�	������u�3��oj��t����P�|,������t����    ����K�F�} u@ǅ\���    j��\���R�E    P�MQ�������u�����U��\����3������M�3��?<����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E���]����U����E�    �} t	�E�   ��E�    �E�E��}� u&hIh�Yj hJ  hHj�P������u̃}� u3�b���    j hJ  hHh,IhI��Z�����   �R  �} t	�E�   ��E�    �U�U�}� u&hlIh�Yj hK  hHj��������u̃}� u3�b���    j hK  hHh,IhlI�jZ�����   ��   � ����u�� ��u�E�   �M�    j j j��URj �E�P� �E��}� u�� P�����3��|h\  h�Ij�M���Q�C�����U��E�8 u3��Q�M�Q�U�Pj��MQj �U�R� ��u,�� P�����j�E�Q�r)�����U�    3���   ��]�����������������������������������������������������������������������������������������������������������������������������U����E�    �} t	�E�   ��E�    �E�E��}� u&h�Ih�Yj h�  hHj��������u̃}� u3�1`���    j h�  hHh�Ih�I�X�����   �X  �} t	�E�   ��E�    �U�U�}� u&hJh�Yj h�  hHj�o������u̃}� u3�_���    j h�  hHh�IhJ�
X�����   ��   �����u�� ��u�E�   �M�    j j j j j��URj �E�P� �E��}� u�� P�����3��~h�  h�Ij�M�Q�������U��E�8 u3��Uj j �M�Q�U�Pj��MQj �U�R� ��u,�� P�O����j�E�Q�'�����U�    3���   ��]���������������������������������������������������������������������������������������������������������������������������������������U����E�Ph�Gj �, ��th H�M�Q�� �E��}� t�UR�U���]�������������������U��EP�7�����MQ�� ]����������������������U����h�P� �E����M��	�U����U��}� t�E��8 tj�M��R�%������j��P�%������    � ��M��	�U����U��}� t�E��8 tj�M��R�[%������j� �P�I%����� �    j���Q�.%����j���R�%�������    ���    �}��t�=h� tj�E�P��$����j�� �h��   k� ��� t+j�   k� ���R�$�����   k� ǁ�    �   �� ��� t+j�   �� ���Q�y$�����   �� ǂ�    �|������Iu'�=|�X�tj�|�R�;$�����|�X���]������������������������������������������������������������������������������������������������������������������������������U����T���EP��>����h�   ����]�����������������U��jjj �B  ��]��������������U��jj j �"  ��]��������������U��Q�= � th ��IU������t�EP� ����!��h�Hh�F�.�����E��}� t�E��Ghq�:����h�Eh @��  ���=T� thT���T������tj jj �T�3���]������������������������������������������������������U��j j�EP�0  ��]������������U��j j j �  ��]��������������U����} t	�E�   ��E�    �E��E��}� u&h��h�Yj h%  hHj�G������u̃}� u3�Y���    j h%  hHh�Hh����Q�����   �   �=� t	�E�   ��E�    �U�U��}� u&h�Hh�Yj h)  hHj��������u̃}� u0�Y���    j h)  hHh�Hh�H�^Q�����   ��M���3���]������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u&h��h�Yj h  hHj��������u̃}� u3�(X���    j h  hHh�Hh���P�����   �   �=� t	�E�   ��E�    �U�U��}� u&h�Hh�Yj h  hHj�c������u̃}� u0�W���    j h  hHh�Hh�H��O�����   ��M���3���]������������������������������������������������������������������������U��Qj � �E��E�P�z,�����M�Q�'�����U�R�p�����E�P�:�����M�Q�C�����U�R�Y�����J����]���������������������������������U��E;Es�M�9 t�U��ЋM���M��]����������U��Q�E�    �E;Es#�}� u�M�9 t
�U��ЉE��M���M�ՋE���]��������������������U��j�����]������������������U��j��H����]������������������U��j�hȅh�Ld�    P���SVW���1E�3�P�E�d�    �[���E�    �=��N  ���   �E����} �  �h�Q� �E��}� ��   �d�R� �E��E�    �E��E؋M�Mк   ����   �E�    �E�    �E���E�M�;M�rj � �U�9u�ދE�;E�s�k�M�R� �E�j � �M��Űh�R� �Eܡd�P� �EԋM�;M�u�U�;U�t�E܉E؋M؉M��UԉUЋEЉE��N���h�Lh�I�������h�Nh�M��������} uj��x3������ t
�+���F���E������   ��} t�,��Ã} t���   �,���MQ�7�����M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������U��j j �EP������]������������U����E�8�t%�M��E��M��U�EB3E��E��M��+���M�Q�E��M��U�EB3E��E��M��+����]������������������������������������U���0�E� �E�   �E���E��M����M�U��B3���E�M�Q�U�R�A������E�H��f�  �U�UЋE�EԋM��UЉQ�E��H�M���U܉U��}����   kE��M�T�U�E�H�M�U��E܃}� ��   �U�M��4���E��E��}� }�E�    �   �   �}� ��   �M�9csm�u)�=� t h��UL������tj�UR�����M����U�M���E��H;M�th���U�R�M����U�� ���E��M܉H�U�R�E�P�)������U�M�I�p(�������&�U��z�th���E�P�M������������E��M���t�U�R�E�P��������E؋�]�����������������������������������������������������������������������������������������������������������������������������U��   ]�������U���H�    ]������������������U���E%�  ���ȋU�����P���E�$�o#����]�����������������U����E��������Dz���]��E�    ��   �E%�  ��   �M����u
�} ��   �E�������]����Au	�E�   ��E�    �U��U��E��u/�M��M�U��   �t	�E���E�M��M�U����U����E%��  f�E�}� t�M�� �  f�Mj ���E�$�"�����]��.j ���E�$�h"�����]��U���  ����-�  �E��M�U���E��]����������������������������������������������������������������������������������U��Q�E%�  ��f�E��M����  f�M��E���]�����������������������U����E�]��E%�  �M���f�E��E���]�������������������������U����E�]�E�  �E��M���  �U����f�M��E��]�����������������������������U��}  �u�} u�   �X�}  ��u�} u�   �B�E%�  =�  u�   �+�M���  ���  u�U����u�} t�   �3�]������������������������������U��Q�E�� t	�E�   �K�M��t	�E�   �:�U��t	�E�   �)�E��t	�E�   ��M��t	�E�   ��E�    �E���]��������������������������S�܃������U�k�l$���   ���3ŉE��C P�KQ�SR�V������u)�E�����E��KQ�SR�CP�KQ�S R�E�P�}�����KQ�'������|����=P� u>��|��� t5�S R���C�$�����$���C�$�CP��|���Q�����$�%���|���R�3����h��  �C P�5�����C�M�3��|$����]��[�����������������������������������������������������������������������������S�܃������U�k�l$���   ���3ŉE��C(P�K Q�SR�������u;�E����E��M������M��C�]��S R�CP�KQ�SR�C(P�M�Q�+�����SR��������|����=P� u?��|��� t6�C(P���C �$���C�$���C�$�KQ��|���R�h����$�%���|���P��1����h��  �K(Q�_4�����C �M�3��)#����]��[��������������������������������������������������������������������������U��Q�E�    �	�E����E��}�}�M��͠�;Uu�E��Ť����3���]������������������U���H�E���E��M��t �U��tj�{<�����E�����E��  �M��t �U��tj�S<�����E�����E��s  �M���   �U���  j�#<�����E%   �E�}�   w�}�   tW�}� t �}�   tv��   �}�   ��   �   �M�������z�p��]���p����]ЋU�E���   �E�������z�p��]��������]ȋM�E���Z�U�������z����]���p����]��E�E���,�M�������z����]��������]��U�E���E�����E��G  �M���;  �U���/  �E�    �E��t�E�   �M���������D��   �U�R�E��� �$�)O�����]؋M��   �M��}�����}�E��x^�]��E�   �   ���]�����Au	�E�   ��E�    �U�U��Eރ�f�E��Mރ�f�M��	�U����U��}����}:�E؃�t�}� u�E�   �M���M؋U܃�t�E�   ��E؋M���M�봃}� t�E����]؋U�E����E�   �}� t
j��9�����E�����E��M��t�U�� tj �9�����E����E��}� t	�E�    ��E�   �E��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��=P� u0�EP���E�$�����$���E�$�MQj�����$�!���E��� !   h��  �UR�z/�����E]������������������������������������U����E�E�]��=P� u1�EP���E��$���E�$���E�$�MQj������$�!��cE��� !   h��  �UR��.�����E���]�������������������������������������U��j �EP�MQ�UR�EP�MQ�UR�0����]����������U���,�E�  ��E�@    �M�A    �U�B    �E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U��t�E��  ��E�H���U�J�E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U���t	�E�    ��E�   �M�����U�B�����M�A�U���t	�E�    ��E�   �M�����U�B�����M�A�U���t	�E�    ��E�   �M������U�B�����M�A�U���t	�E�    ��E�   �M܃���U�B�����M�A�U��� t	�E�    ��E�   �M؃��U�B�����M�A�z0���E��U���t�E�H���U�J�E���t�M�Q���E�P�M���t�U�B���M�A�U���t�E�H���U�J�E��� t�M�Q���E�P�M���   �U�}�   w�}�   t+�}� tI�}�   t.�K�}�   t�@�E����U�
�1�E�������U�
��E�������U�
��E�����U�
�E���   �M�t5�}�   t�}�   t�1�U����M��"�U������M���U������M��U���  ���E��� ��ʋU�
�}  tT�E�H ���U�J �E�H ���U�J �E�M��X�U�B`���M�A`�U�B`���M�A`�U�E� �ZP�X�M�Q ���E�P �M�Q �����E�P �M�U��Y�E�H`���U�J`�E�H`�����U�J`�E�M��XP�B���URjj �E�P�8 �M�Q����t�E�����U�
�E�H����t�U�����M��U�B����t�M�����E��M�Q���t�E����U�
�E�H��t�U���ߋM��U����Eԃ}�w[�M��$�T,�U�%����   �M��;�U�%����   �M��%�U�%����   �M���U�%�����M��U������E�t�}�t �}�t2�@�M���������   �E��(�M���������   �E���M��������E��}  t�M�U�BP���E�M�AP���]Ð�+�+�+�+����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�EP�MQ�UR�EP�MQ�UR��(����]����������U��Q�E�E��}�t�}�~ �}�~��=��� !   ��=��� "   ��]�����������������������U��� �EP�!������E�}� t^�M�M��U�U�E�E�M�M��U�U�E �E��M$�M�h��  �U(R��&�����E�P�z������u�MQ�$�����E��"� h��  �U(R�&�����EP��#�����E ��]����������������������������������������������������U��Q�= �|����E��E���?�E������E�    �E���]��������������U����= �|8�i���E��E#E�M��#M���E��U������U��U��E�P�'�������E�    �E���]����������������������������U��Q�= �|�]��e���U���]��������������������U��Q�= �|�]���E�    �E���]����������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �e�= ���   �E��@tp�=Ъ tg�E�    �U�E������Q�M���E�}�  �t�}�  �t	�E�    ��E�   �E�Ëe��Ъ    �M�ΈM�U�E�������U�⿉U�U�M�d�    Y_^[��]����������������������������������������������������������U��Q����E��E��?E��E��M�Q�h�������]�������������������������U��Q�= �|�K���E��E���?�E���E�    �E���]�������������������U��Q�}����E���]����������������U�����}��E#E�M��U��#��f�E��m��E���]���������������������U����E��t
�-���]���M��t����-���]������U��t
�-Ī�]���E��t	�������؛�M�� t���]����]����������������������������U��Q��}��E���]�����������������U���0���3ŉE�SV� �    �ܪ���ܪj
��
�����[  �E�    �E�    �E�    � �   �ܪ���ܪ�u�3�3����^�N�V�   k� �L��Mк   �� �D�5Genu�   k��L���ineI��   ��L���ntel�u	�E�   ��E�    �UԈUߍu�   3����^�N�V�   k��   k� �L��L�   ��   �� �L��L�   k� �L��M��U߅�to�E�%�?�=� tS�M؁��?���` tB�U؁��?���p t1�E�%�?�=P t"�M؁��?���` t�U؁��?���p u�$����$��}�|O�u�   3����^�N�V�   �� �   ��D��D�   �� �T���   t�$����$��   �� �T���   ��   � �   �ܪ���ܪ�   �� �T���   tV�   �� �L���   tB� �   �ܪ���ܪ�   ���L��� t� �   �ܪ�� �ܪ3�^[�M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������̅�uf���fn�f`�fa�fp� SQ�ك���ux�ڃ���t0ffAfA fA0fA@fAPfA`fAp���   KuЅ�t7����t��I f�IKu���t����t
f~�IJu���t�AKu�X[��ۃ�+�R�Ӄ�t�AJu���t
f~�IKu�Z�^�����������������������������������������������������������U���0�} t�} v	�E�   ��E�    �E�E��}� u#hKh�Yj jhxKj�4�������u̃}� u0�u4���    j jhxKh�KhK��,�����   �k  �} ��   �U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U�E�Ph�   �M��Q������} t	�E�   ��E�    �U�U�}� u#h�Kh�Yj jhxKj�Z�������u̃}� u0�3���    j jhxKh�Kh�K��+�����   �  �M�M��U�U��E��M���E���MЋU����U��E���E�}� t�M����M�t�ȃ}� ��   �U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U��E�Ph�   �M��Q������ L��t3�t	�E�   ��E�    �M܉M؃}� u#hPLh�Yj jhxKj�5�������u̃}� u-�v2��� "   j jhxKh�KhPL��*�����"   �o�}�tg�}���t^�E+E���;EsP�M+M����U+�9h�s
�h��E���M+M����U+щUԋE�Ph�   �M+M��U�D
P�����3���]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u#h �h�Yj j)h�Lj�z�������u̃}� u+�0���    j j)h�Lh�Lh ��)���������U�B��]�������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u�����     �0��� 	   �����  �} |�E;<�s	�E�   ��E�    �M��M܃}� u#hMh�Yj j.h�Mj�j�������u̃}� u9�����     �/��� 	   j j.h�Mh�MhM��'��������9  �E���M������0��D
��t	�E�   ��E�    �M؉Mԃ}� u#h�Mh�Yj j/h�Mj���������u̃}� u9�����     �/��� 	   j j/h�Mh�Mh�M�_'��������   �EP�3�����E�    �M���U������0��L��t�UR�0�����E��9�.��� 	   �E�����3�u#h(Nh�Yj j9h�Mj��������u��E������   ��UR������ËE�M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������U��QV�EP���������tn�}u�   k� ��0����   ��u�}u1�   k� ��0��QD��tj��������j������;�t�EP������P�� ��t	�E�    �	�� �E��MQ�������U���E������0��D �}� t�U�R�D���������3�^��]����������������������������������������������������������������������U��} u#h�Nh�Yj j.h Oj���������u̋M�Q��   tK�E�H��t@j�U�BP�j������M�Q�������E�P�M�    �U�B    �E�@    ]������������������������������������������U��j�h(�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u�+��� 	   �����  �} |�E;<�s	�E�   ��E�    �M��M܃}� u#hhOh�Yj j,h�Oj���������u̃}� u.�+��� 	   j j,h�OhPPhhO�s#��������X  �E���M������0��D
��t	�E�   ��E�    �M؉Mԃ}� u#hdPh�Yj j-h�Oj�B�������u̃}� u.�*��� 	   j j-h�OhPPhdP��"���������   �EP�3/�����E�    �M���U������0��L��t;�UR������P�� ��u�� �E���E�    �}� u�C������M���)��� 	   �E�����3�u#h(Nh�Yj jEh�Oj�g�������u��E������   ��MQ������ËE�M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������U��j�hH�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u�����     �(��� 	   �����  �} |�E;<�s	�E�   ��E�    �M��M܃}� u#hMh�Yj jBh�Pj���������u̃}� u9�6����     �0(��� 	   j jBh�PhQhM� ��������L  �E���M������0��D
��t	�E�   ��E�    �M؉Mԃ}� u#h�Mh�Yj jCh�Pj�\�������u̃}� u9�����     �'��� 	   j jCh�PhQh�M����������   �EP�B,�����E�    �M���U������0��L��t�UR�EP�MQ�������E��D�'��� 	   �����     �E�����3�u#h(Nh�Yj jNh�Pj��������u��E������   ��MQ�8�����ËE�M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������U�츔<  �,�����3ŉE�ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    �} u3��C  �} tǅ|���   �
ǅ|���    ��|��������������� u#hQh�Yj jlh�Pj��������u̃����� u9�T����     �N%���    j jlh�Ph<QhQ���������  �U���E������0��T$������������������t����������   �U��uǅ����   �
ǅ����    ��������x�����x��� u#h`Qh�Yj jth�Pj�C�������u̃�x��� u9�|����     �v$���    j jth�Ph<Qh`Q�����������  �U���E������0��T�� tjj j �EP������MQ���������   �U���E������0��T��   tt������p�����p����Hl�   �⃼�    uǅ����   �
ǅ����    ��������������l���Q�U���E������0��R�� ������������ �  ������ t����������  �� ��t���3�f������ǅ����    ǅ����    �U������������+E;E��  ǅ����    ���������  ���������
uǅ����   �
ǅ����    �������������U���E������0��|8 ��   �U���E������0��T4R�%������u&h�Qh�Yj h�   h�Pj��������u̋M���U������0��   k� �T4�T��   �� ��������T�E���M������0��D
8    j�E�P������Q�� �������u�{  ��   �������P�%��������   ������+M�U+у�v3j������P������Q�v �������u�'  ���������������T�E���M������0�������� �D
4�M���U������0��D8   ����������������  �"j������R������P����������u�  ���������������e��������t��������uM������f�f��������������
uǅ����   �
ǅ����    �����������������������������������P  j j j�M�Qj������Rj ��t���P� ������������ u��  �sj ������Q������R�E�P�M���U������0��Q�� ��t*������+U�����������������;�����}�  ��� �������n  ������ ��   ǅ����   �   k� �D�j ������P������Q�U�R�E���M������0��
P�� ��t3������;�����}��   ������������������������������� ��������   ��   ��������t����������   ������P�������������;�u����������������� �������p������ tbǅ����   �   f������������R�)������������;�u ������������������������������� ��������D����7  �M���U������0��L��   ��  ǅ����    ���������[  ǅ����    ǅ����    �E������������+M;M�'  ������������������������+�=�  ��   ������+U;Usr�����������������������������������
u'���������������������������������������������������������������g���j ������Q������������+�R������Q�U���E������0��R�� ��t,�����������������������������+�9�����}���� �������������A  ���������[  �M������ǅ����    ������+U;U�1  ������������������������+ʁ��  ��   ������+E;Es{������f�f����������������������������
u,���������������   ������f���������������������f������f����������������]���j ������P������������+�Q������P�M���U������0��Q�� ��t,�����������������������������+�9�����}���� �������������  �U������ǅ����    �E������������+M;M��  ǅ����    ��H�����������������H���+�=�  sz������+U;Usl������f�f����������������������������
u�   ������f�
��������������������f������f����������������q���j j hU  ������Q��������H���++���P��H���Pj h��  � ������������ u�� �������   �   ǅ����    j ������Q������+�����R������������Q�U���E������0��R�� ��t�������������������� �������������;������������;�����~�������+E�������F����Yj ������Q�UR�EP�M���U������0��Q�� ��tǅ����    ��������������� ������������ ��   ������ t9������u����� 	   �������������������R�[���������\�L�E���M������0��D
��@t�M���u3��+�����    �����     �����������+������M�3��������]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���V�E�    �} t	�E�   ��E�    �E��E�}� u#ht�h�Yj jmh�Qj�b�������u̃}� u.����    j jmh�Qh4Rht�� ���������  �U�U��E��H��   t�U��B��@t����  �M��Q��t�E��H�� �U��J����  �E��H���U��J�E��H��  u�U�R�w������E��M��Q��E��HQ�U��BP�M�Q�����P��������U��B�E��x t	�M��y�u:�U��z t	�E�    ��E�   �E��HM��U��J�E��@    �����   �M��Q��   u�E�P� �������t@�M�Q� �������t/�U�R�o ���������E�P�^ ���������0��E���E���M��Q��   ���   u�E��H��    �U��J�E��x   u#�M��Q��t�E��H��   u
�U��B   �E��H���U��J�E������   �U�E�����U��
�E�^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hh�h�Ld�    P�ĄSVW���1E�3�P�E�d�    j�Z������E�    h�   hHRjj@j �������E�}� u"�E�����j��E�Ph���M�����E��G  �   k� �E䉂0��<�    �	�M��@�M�   k� ��0���   9M�su�U��B �E�� �����M��A
�U��B    �E�H$�ဋU�J$�E�H$���U�J$�   k� �U��D
%
�   �� �M��D%
�U��B8    �E��@4 �i�����t���Q�� �U�����  �}� ��  �E���M܋U����UԋE�E܉E؁}�   }�M܉M���E�   �UĉU��E�   �	�EЃ��EЋ<�;M���   h�   hHRjj@j �G������E�}� u�<��U��   �EЋM��0��<��� �<��	�E��@�E�MЋ�0���   9U�sf�E��@ �M�������U��B
�E��@    �M�Q$�​E�P$�   k� �E��D%
�   �� �U��D
%
�E��@8    �M��A4 �|��������E�    ��U����U��Eԃ��EԋM؃��M؋U�;U���   �E؃8���   �M؃9�ty�U����tn�M����u�E؋Q�� ��tS�U����E������0��E�M�U؋��M�UԊ�Aj h�  �M��Q��������U�B���M�A�G����E�    �	�U����U��}��H  �   k� �U����0��U�E�8�t�M�9��  �U��B��}� u	�E�������}�u	�E�������E������E��E��M�Q�� �Ẽ}����   �}� t�U�R�� �Eȃ}� tl�E�M̉�Uȁ��   ��u�E��H��@�U�J��E�%�   ��u�M��Q���E�Pj h�  �M��Q��������U�B���M�A�5�U��B��@�M�A�U�������=|� t�E��|����B������E��H�ɀ   �U�J�����E������   �j�/ �����3��M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    �	�E����E��}�@}y�M��<�0� tg�U���0��E��	�M���@�M��U���0�   9E�s�M��y t�U���R� ��j�E���0�Q�������U���0�    �x�����]������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�   ��E�    �E�E��}� u#h �h�Yj j0hxRj�2�������u̃}� u.�s
���    j j0hxRh�Rh ��������������F�UR�B������E�    �EP�������E؉U��E������   ��MQ�� ����ËE؋U܋M�d�    Y_^[��]����������������������������������������������������������������������������������U��\  ������3ŉE�V�} u#ht�h�Yj jZhxRj��������u̋M������������R�m������������������x }�������A    jj j ������R������������������������� |	������ s�������[  ��������������������0��D
$�����������������Q��  u#�������@�������+ȋ�����������  �������������
+H�������������B���  ����������  ��������������������0��|0 �m  �������������
+H�鉍�����������z u�������������g  �2  j ��������������������0��D
,P�L
(Q������R��������������������������������������0�������������������������������;T(u������������������;T,t�������  j ������Ph   ������Q��������������������0��R�� ��u�������r  j ������P������Q������R������������������������ |	������ s�������(  ������;�����v�������  �������������������������������������������� ��   ������������9�����ss���������u5������������9�����s�������Q��
u������������������������X���������������������������P���������������+Ћ�3������������0  ��������������������0��L��   tO�������B���������������������������������;s���������
u�����������������'�������Q��   u�.���    �������  �����������u3ҋ������t  �������Q���4  �������x uǅ����    �  �������������+B������A��������������������������0��T��   ��  jj j ������P�F�����������������������;�������   ������;�������   �������H������������������B���������������������������;�����s���������
u���������������ċ������H��    t����������������   j ������P������Q������R�p����������������������� |	������ s��������   ������   w*�������H��t�������B%   uǅ����   ��������Q��������������������������0��D
��t����������������������u�������艅����3ɋ�����+��������������������������������u�������ꉕ����������3�����������^�M�3��������]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} u#ht�h�Yj jdh�Rj�6�������u̋M�M��U�R�������E��E��H��   u$�Z ��� 	   �U��B�� �M��A����X  �-�U��B��@t"�+ ��� "   �M��Q�� �E��P����)  �M��Q��tH�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J�����  �E��H���U��J�E��H���U��J�E��@    �E�    �M�M��U��B%  uC�
����    �� �9E�t������    ���9E�u�E�P���������u�M�Q�������U��B%  ��   �M��U��+By&h`Sh�Yj h�   h�Rj覸������u̋U��E��
+H�M�U��B���M���U��B���M��A�}� ~�U�R�E��HQ�U�R��������E��q�}��t!�}��t�E����M������0��M���E���U��B�� t7jj j �M�Q�,������E�U�U�#U���u�E��H�� �U��J����O�E��H�U���E�   �E�P�MQ�U�R�N������E��E�;E�t�M��Q�� �E��P�����E%�   ��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E������E������}�u!�ӻ���     ������ 	   ��������  �} |�E;<�s	�E�   ��E�    �M�M��}� u#hMh�Yj j@h�Sj� �������u̃}� u<�\����     �V���� 	   j j@h�Sh\ThM�������������`  �E���M������0��D
��t	�E�   ��E�    �M܉M؃}� u#h�Mh�Yj jAh�Sj��������u̃}� u<軺���     ����� 	   j jAh�Sh\Th�M�������������   �EP�b �����E�    �M���U������0��L��t �UR�EP�MQ�UR�)������EЉU��K�1���� 	   �!����     �E������E�����3�u#h(Nh�Yj jLh�Sj蟴������u��E������   ��UR�J�����ËEЋUԋM�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EP芽�����E��}��u:������ 	   3�u#h(Nh�Yj jwh�Sj�x�������u̃������s�EP�M�Q�UR�EP�M�Q�� ��u�� P�������������>�U���E������0��T����E���M������0��T�E�U���]�����������������������������������������������������U����} u#ht�h�Yj j.hxTj薲������u̋\����\��U�U�j:h�Tjh   臮�����E��E��M��H�}� t�U��B���M��A�U��B   �%�E��H���U��J�E����M��A�U��B   �E��M��Q��E��@    ��]������������������������������������������������������������U��j�hȆh�Ld�    P���SVW���1E�3�P�E�d�    �E�    j�s������E�    �E�   �	�E���E�M�;����   �U�|��<� t|�M�|����H��   t"�U�|���Q�f��������t	�U����U��}�|=�E�|����� R� j�E�|���R�}������E�|���    �Y����E������   �j������ËE��M�d�    Y_^[��]���������������������������������������������������������������������������U���0�} t�} v	�E�   ��E�    �E�E��}� u#hUh�Yj jhxKj��������u̃}� u0�E����    j jhxKhtUhU�������   �w  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R�z������} t	�E�   ��E�    �E�E�}� u#h�Kh�Yj jhxKj�&�������u̃}� u0�g����    j jhxKhtUh�K��������   �  �U�U��E�E��M��Uf�f��M���UЋE����E��M���M�}� t�U����U�t�ƃ}� ��   3��Mf��}�tJ�}���tA�}v;�U��9h�s
�h��E��	�M���M��U���Rh�   �E��P�W������ L��t3�t	�E�   ��E�    �E܉E؃}� u#hPLh�Yj jhxKj���������u̃}� u-�=���� "   j jhxKhtUhPL�������"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9h�s�h��U���E+E����M+ȉMԋU���Rh�   �E+E��M�TAR�h�����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�E��M�Q�UR�EP�MQ��������]�����������U��Q�E�E��M�Q�UR�&�������]�������������������U��Q�E�E��M�Q�UR�EP肭������]���������������U��Q�E�E��M�Q�UR�`�������]�������������������U��Q�E�E��M�Q�UR�EP�g�������]���������������U��Q�E�E��M�Qj �UR�EP�MQ�UR��������]���������������������U��Q�E�E��M�Q�UR�EP�MQ�UR�EP�=�������]�������������������U���L�E�    3��E��E��E��EĉEȉẺEЍM��M��} t	�E�   ��E�    �U��U�}� u&h��h�Yj h�   h�Uj裪������u̃}� u1������    j h�   h�Uh�Uh���>���������o  �} t	�E�   ��E�    �M��M�}� u&hX�h�Yj h�   h�Uj�$�������u̃}� u1�e����    j h�   h�Uh�UhX������������   �E�E܋M��AB   �U��E�B�M��U��E��@����M�Qj �UR�E�P��������E��} u�E��   �M��Q���U�E��M�H�}� |"�U���  3Ɂ��   �M؋U�����M����U�Rj �������E؋E��H���M�U��E�B�}� |!�M��� 3�%�   �EԋM�����E����M�Qj �J������EԋE���]�����������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�E��M�Qj �UR�EP�MQ���������]�������������������������U��Q�E�E��M�Q�UR�EP�MQ�UR踱������]�����������������������U��Q�E�E��M�Q�UR�EP�MQ�UR��������]�����������������������U��Q�E�E��M�Qj �UR�EP�MQ�خ������]�������������������������U��������d]����U��l�P� ]����������������U���t�����`]����U��E�d��M�h��U�l��E�p�]����������U��j�h(�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    j 蜧�����E�    �} u�E�d��E��Q� �E��E�   ��E�h��U��P� �E��E�   �}� t�}�tj � �M���E������   �j ������Ã}� u3���}�t
�U�R�U���   �M�d�    Y_^[��]� ��������������������������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�    �E�    �E�    �E�    �E�EԋMԃ��Mԃ}���   �U�����$�܂�E�d��M��U��E؃��E��  �E�h��M��U��E؃��E���   �E�l��M��U��E؃��E���   �E�p��M��U��E؃��E��   �����E܃}� u�����  �M܋Q\R�EP��  �����E�M��U��   �}3�t	�E�   ��E�    �M̉Mȃ}� u&h<Vh�Yj h�  h�Vj�9�������u̃}� u1�z����    j h�  h�Vh�Vh<V�����������5  �E�P� �E��}�u3��  �}� uj�ڥ���}� t
j 躤�����E�    �}t�}t�}u,�M܋Q`�UċE��@`    �}u�M܋Qd�U��E��@d�   �}u:�Hz�M��	�UЃ��UСHzLz9E�}kM��U܋B\�D    ���j � �M��E������   ��}� t
j �m�����Ã}u�U܋BdPj�U����
�MQ�U����}t�}t�}u�U܋EĉB`�}u	�M܋U��Qd3��M�d�    Y_^[��]Ë�d�؀������� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�E��M��Q;Ut�E����E�k@zM9M�s��k@zU9U�s�E��H;Mu�E���3���]���������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�    �}t�}u�R  �}t�}t�}t�}t
�}�F  j 財�����E�    �}t�}u=�=t� u4jh�~�� ��u�t�   ��� ���å���0�E�   �E�E؋M؃��M؃}���   �U���ȇ�$����d�Q� �E܃}t�UR� �d��r�h�P� �E܃}t�MQ� �h��L�l�R� �E܃}t�EP� �l��%�p�Q� �E܃}t�UR� �p��E������   �j �������Ã}� t��   ��   �}t�}t�}t��   ������E��}� u��   �E��x\�yuLhZ  hVj�DzQ�R������E̋U��ẺB\�}� t�DzQh�y�U��B\P�J�������h�M��Q\R�EP�@������E�}� u�J�M�Q�U܃}t3�E�H;Mu(�U�E�B�M���M�k@z�E�P\9U�r��͋E��   �M�MԋUԃ��Uԃ}�w�E�����$�������}3�t	�E�   ��E�    �EȉEă}� u&h<Vh�Yj h�  h�Vj�,�������u̃}� u.�m����    j h�  h�Vh�Vh<V���������������M�d�    Y_^[��]Ë�L�����s�� �I �#�     �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���`���3ŉE��E�    j � �E��E�    �E�    �����E��E�    �=�� ��   h   j hW�� �E�}� u�� ��Wuj j hW�� �E�}� u3��q  h$W�E�P�� �E�}� u3��R  �M�Q� ���h4W�U�R�� P� ���hHW�E�P�� P� �|�h`W�M�Q�� �E�U�R� ����=�� th�W�E�P�� P� ����  ��t �} t
�MQ�� �}� t
�   �  �}� ��   ���R� �E��E�    �E��E��M�M��U�U��E�E�3ɉM��}� u3��S  j j �U�Rh�*j j �� �E؃}� u3��,  j j��E�P�� ��u�E��  3��  ���;M�th���;U�t]���P� �Eԋ��Q� �E��}� t8�}� t2�UԉE܃}� t�U�Rj�E�Pj�M�Q�U���t�U���u�E�   �}� t�E    �E�W���;M�t���R� �E��}� t�U��E�}� t*�|�;E�t �|�Q� �EЃ}� t
�U�R�UЉE䡈�P� �Eȃ}� t�MQ�UR�EP�M�Q�U���3��M�3��]�����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�E��M��QR�E��HQ�U��BPj �M���ҋM��A3���]� ��������������������������U���]�����������U��8�]�������U����} |�}}	�E�   ��E�    �E��E��}� u*h�Wh�Yj h�   h Xj��������u�����}� u0�>����    j h�   h Xh�Yh�W������������c�}�u�U��8��Q�E��8��M�}�uj��� �U��8��'�}�uj��� �M��8���U�E��8��E��]����������������������������������������������������������������������������U��Q�8��E��M�8��E���]���������������������U����} |�}}	�E�   ��E�    �E��E��}� u'h�Wh�Yj jsh Xj蔖������u译���}� u.������    j jsh Xh`Xh�W�.���������   �}�t�U���t	�E�    ��E�   �E�E��}� u'h�Xh�Yj jxh Xj��������u�*����}� u+�L����    j jxh Xh`Xh�X����������/�}�u�U��,���E��,��M�U�E��,��E��]�����������������������������������������������������������������������������������U��j�hH�h�Ld�    P���LP  �	������1E�3ŉE�SVWP�E�d�    ǅܯ��    ǅ���    ƅ���� h�  j ������P�������ƅ���� h�  j ������Q�ٻ����3�f�����h�  j �����P躻����ƅ���� h�  j ������Q蝻�����} |�}|����t  �E�    �}��   �D��   ��@����   j h  h Xh�Yh�Yj
h   ������Q�UR�w�����P������hPZ�� �} t�E�������
ǅ�����Z������Q�� h�Z�� ������R�� h�4�� �ݎ��ǅܯ�������  �} ��   ǅ̯��    ������ ������������     �M Q�URh�  h   ������P��������̯����̯�� }*j h-  h Xh�Yh��j"j�����Q虐���� �p������������̯�� }8j h0  h Xh�Yh�ZhX[h   ������P�i�����P觝�����}uV�} tǅ����\\�
ǅ����t\j h5  h Xh�Yh�[������Qh   ������R������P�K�����j h7  h Xh�Yh�\������Ph   ������Q�F�����P�������}u�U��,���t8j h<  h Xh�Yh ]hX]h   ������Q�������P�Ĝ����j h=  h Xh�Yh`]h�4h   ������R�������P茜�����} ��   ǅЯ��    ������ ������������     ������Q�UR�EPh�]h�  h   ������Q��������Я����Я�� }*j hD  h Xh�Yh��j"j�����R螎���� �u������������Я�� }8j hG  h Xh�Yh�]hX[h   ������R�n�����P講�����:j hK  h Xh�Yh�^������Ph   ������Q�2�����P�p�����ǅ����    ǅȯ��    j�������Rh   �����P������Q��������ȯ��j hP  h Xh�Yh�^j"j��ȯ��R譍���� ��ȯ�� t8j hR  h Xh�Yh�_h�`h   �����P�+�����P�Ț�����=4� u�=$� �#  ǅԯ��    ǅد��    j跐�����E�   �4���ԯ�����ԯ���B��ԯ����ԯ�� tHǅ����    ������Q������R�EP��ԯ���Q�҃���tǅ���   ��������ܯ���렃���� un�$���د�����د���B��د����د�� tHǅį��    ��į��Q�����R�EP��د���Q�҃���tǅ���   ��į����ܯ�����E�    �   �j������Ã���� ��  �=8� t?ǅ����    ������Q������R�EP�8�����tǅ���   ��������ܯ������� �4  �U��,���t>�M�<�8��t1j ������R������P�W�����P������Q�U��8�P�� �M��,���t������P�� �M��,�����   �   k� ������������   s�����������Ƅ���� �} t9j h�  h Xh�Yh�Yj
h   ������P�MQ�������P�C������} t�������������
ǅ����    ������P�MQ������R�EP�MQ�UR��������ܯ���E������   ��}u�D������Ë�ܯ���M�d�    Y_^[�M�3�貫����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hx�h�Ld�    P���T�  �y������1E�3ŉE�SVWP�E�d�    ǅ���    ǅ���    3�f������h�  j ������Q�d�����3�f�����h�  j �����P�E�����ƅ���� h�  j ������Q�(�����3�f�����h�  j �����P�	������} |�}|����v  �E�    �}��   �D��   ��B����   j h�  h Xhah@aj
h   ������P�MQ�b�����P�Q�����h�a�� �} t�U������
ǅ����a�����P�� h b�� ������Q�� h4b�� �I���ǅ��������  �} ��   �X����������K����     �E P�MQh�  h   �����R�a��������������� }*j h  h Xhah��j"j������ P������ ���������������� }8j h
  h Xhah8bh��h   �����R������P�������}uV�} tǅ����c�
ǅ����cj h  h Xhah�b�����Ph   ������Q�$�����P�������j h  h Xhah d�����Rh   ������P�������P臒�����}u�M��,���t8j h  h Xhah�dh�dh   ������P�t�����P�:�����j h  h Xhah�dh4bh   ������Q�<�����P�������} ��   ǅ���    �i����������\����     ������P�MQ�URhHeh   h   �����P誩�������������� }*j h   h Xhah��j"j������Q������ ���������������� }8j h"  h Xhah�h��h   �����P������P�"������:j h&  h Xhahhe������Qh   �����R�I�����P������ǅ���    j h,  h Xhah�ej"jj������Ph   ������Qj 辢����P�>����� ���������� t8j h.  h Xhah�fhpgh   ������R������P�S������=4� u�=$� �!  ǅ���    ǅ���    j�B������E�   �4�������������Q���������� tHǅ���    �����P������Q�UR������H�у���t����������ǅ���   �렃���� um�$�������������Q���������� tHǅ���    �����P�����Q�UR������H�у���t����������ǅ���   ���E�    �   �j製����Ã���� ��  �=8� t?ǅ���    �����P������Q�UR�8�����t����������ǅ���   ����� �W  �M��,����[  �E�<�8���J  �M��8�R�� ����������t�Jj �����P�����Q�B�����P�����R�E��8�Q�� ��t��   �� ��t��   ǅ���    j h�  h Xhah�gj"jj������Rh   �����P�����Q�������P�}����� ���������� t>�����Pt5j �����R�����P菬������P�����Q�U��8�P�� �@����� v������������j �����R�����P�����Q�U��8�P�� �M��,���t�����P�� �M��,�����   �   k� ����������    s������3ҋ����f�������} t9j h�  h Xhah@aj
h   ������Q�UR辻����P譌�����} t������������
ǅ���    �����Q�UR�����P�MQ�UR�EP�Y�����������E������   ��}u�D������Ë�����M�d�    Y_^[�M�3�������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � �����������������������U��Q�E�   ���U�zx t�E�Hx�   ���E���    t�M���   �   ���M�y| t�U�B|�   ���U���    t�E���   �   ���E�    �	�E����E��}�q�M����U�|
��t&�E����M�| t�U����E�L�   ���E����M�| t&�U����E�| t�M����U�D
�   ��뀋U���   �   �   ����]���������������������������������������������������������������������������������U��Q�E���    ��   �M���   (���   �U�zx ��   �E�Hx�9 ��   �U���    t4�E���   �9 u&j�U���   P�o������M���   R�l������E�x| t.�M�Q|�: u#j�E�H|Q�8������U���   P������j�M�QxR������j�E���   Q�������U���    to�E���   �9 uaj�U���   -�   P�Ί����j�M���   ��   R贊����j�E���   ��   Q蚊����j�U���   P膊�����M���   ��t8�U���   ���    u&�M���   R�w�����j�E���   Q�?������E�    �	�U����U��}��  �E����M�|��tR�U����E�| tB�M����U�D
�8 u0j�M����U�D
P�։����j�M��U����   P辉�����M����U�|
 t�E����M�| uF�U����E�| u�M����U�|
 t&h`hh�Yj h�   hPjj�z������u̋M����U�|
 t:�E����M�| t*�U����E�L�9 uj�U����E�LQ�����������j�UR���������]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�} �  �E������U�zx t�E�Hx������E���    t�M���   ������M�y| t�U�B|������U���    t�E���   ������E�    �	�E����E��}�m�M����U�|
��t$�E����M�| t�U����E�L������E����M�| t$�U����E�| t�M����U�D
�����넋U���   �   ������E��]������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �0����E��E��Hp# �t	�U��zl uDj�x�����E�    �4�P�M���lQ�B������E��E������   �j���������ͩ���Pl�U�}� u
j �#������E�M�d�    Y_^[��]�������������������������������������������������������U��Q�} t�} u3��\�E��M��U�;UtI�E�M��UR�������}� t�E�P�������}� t�M��9 u�}�8�t�U�R��������E��]���������������������������������������������U��=l� uj�艒�����l�   3�]�������������U��Q�E�E��M���  �M��}�wP�U���ȯ�$����   k� ���j�1�   �� ���j�!�   �዁�j��   k����j�3���]Ë�m�}������� �����������������������������������������������������U��j�h�d�    P��$���3�P�E�d�    �E�    �E�P�M�����E�    ���    �}�u)���   ��E��E������M������E��}�c�}�u)���   ��E��E������M������E��N�4�}�u.���   �M��������Q�U��E������M�蹎���E���E�E��E������M�蟎���E��M�d�    Y��]�������������������������������������������������������������������������������U��Q�E�    �	�E����E��}�  }�MM��A ��U�B    �E�@    �Mǁ      �E�    �	�U����U��}�}3��M��Uf�DJ���E�    �	�E����E��}�  }�MM��U���p��A���E�    �	�M����M��}�   }�UU��E���q���  �׋�]���������������������������������������������������������U���   ���3ŉE�������P�M�QR�L ���J  ǅ����    ���������������������   s�������������������и   k� Ƅ���� �   k� ������������������������������������tP�����������������������������������B9�����w������   s������Ƅ���� ���j �U�BP������Qh   ������Rjj �˩����j �E�HQh   ������Rh   ������Ph   �M��  Rj 質����$j �E�HQh   ������Rh   ������Ph   �M��  Rj �y�����$ǅ����    ���������������������   ��   ��������M������t:�E������H���U������J�E�������������������  �]��������E������t:�U������B�� �M������A�U�������������������  ��U�����Ƃ   �2�����   ǅ����    ���������������������   ��   ������Ar?������Zw6�M������Q���E������P�������� �U�������  �X������ar?������zw6�E������H�� �U������J�������� �M�������  ��U�����Ƃ   �<����M�3�薎����]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hȇh�Ld�    P���SVW���1E�3�P�E�d�    �E�    � ����E��E��Hp# �t�U��zl ��   j�o�����E�    �E��Hh�M�U�;|�tK�}� t$�E�����Iu�}�X�tj�U�R��|�����E��|��Hh�|��U�E�   ���E������   �j�e�������	�U��Bh�E�}� u
j 誂�����E�M�d�    Y_^[��]������������������������������������������������������������������������������U����E�    �E�P�M��<w���M�肺���H�y t �M��q����P�B�E��M��\����E����E�    �M��F����E���M��9�����]���������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E����������E�������E܋Hh�M��UR�*������E�E��M;H�  h[  h�jjh   �h�����E��}� ��  �Uܹ�   �rh�}��E��     �M�Q�UR�m�����E؃}� ��  �E܋Hh�����Ju�E܁xhX�tj�M܋QhR�z�����E܋M��Hh�U܋Bh�   ���U܋Bp���1  � ����"  j��l�����E�    �U��B����M��Q����E���  ����E�    �	�U���U�}�}�E�M�U�f�LJf�E�����E�    �	�U���U�}�  }�E�E�M�P��P����E�    �	�E���E�}�   }�M�M�U䊁  ��X��׋|������Ju�=|�X�tj�|�P�y�����M��|��U�   ���E������   �j��������(�}��u"�}�X�tj�M�Q�5y���������    ��E�    �E؋M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���,���3ŉE�V�EP�&������E�} u�MQ�a�����3��0  �E�    �	�Uԃ��Uԃ}��t  kE�0����;M�\  �E�    �	�U���U�}�  s�EE��@ ���E�    �	�M����M��}���   kU�0�E�����M��	�U܃��Uܸ   k� �U��
��ts�   �� �U��
��t`�   k� �E���M��	�U���U�   �� �M��9U�w*�}�   s!�E���x��UU��B��MM�A��q����F����U�E�B�M�A   �U�BP��������M��  �E�    �	�U����U��}�skE�0�M��U�u�f��p��f�DJ�ՋMQ�������3��  �y����} t!�}��  t�}��  t�UR� ��u����q  �E�P�MQ�L ���?  �E�    �	�U���U�}�  s�EE��@ ��M�U�Q�Eǀ      �}���   �M�M��	�U؃��U؋E����tE�U��B��t:�M���U��	�E���E�M��Q9U�w�EE��H���UU�J����E�   �	�E���E�}��   s�MM��Q���EE�P�֋M�QR�|������M��  �U�B   �
�E�@    �E�    �	�M����M��}�s3ҋE��Mf�TA��UR�Z�����3���=�� t�EP�1�����3�����^�M�3�������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��}�|	�}�   ~#h�jh�Yj j8h0kj�0e������u̋MQ�URj �a����]������������������������U����EP�M��n���}�|	�}�   ~#h�jh�Yj jDh0kj��d������u̃}�|5�}�   ,�M�踱������   �M�H#U�U��M��~���E��9�/�M�茱��� �   k�����   �#M�M��M��f~���E���M��Y~����]�������������������������������������������������������U��=� u�E�ȳ�A#E��j �UR�EP��w����]�����������������������������U���0�EP�M��sm���}�|6�}�   -�M�誰������   �E�B#M�M�M��}���E���   �M��}���P�U�����   R臱������tN�E��%�   �   k� �D��   �� �M�L��   ��U�}�s������E��D� �E�   �2�   k� �E�D��E�   �}�s�谡���M��D� �E�   j�M��ٯ����BP�M�Q�U�R�E�Pj�M�软��P�r�������u�E�    �M��|���E���M�#M�M��M��|���E���]�������������������������������������������������������������������������������������������������U��QV�E�    �} u�4�EPj ���Q��E��}� u�� P�ړ�����������0^��]��������������������U���V�E�E��} u�MQ��������   �} u�UR�'�����3��   �E�    �}�w)�} u�E   �EP�MQj ���R��E���EP趙�����}����    3��e�}� u	�=�� u%�}� t��� P���������F����0�E��1�MQ�g�������u�� P�ؒ�����������03���J���^��]�������������������������������������������������������������������������U���V�} t	�E�   ��E�    �E��E�}� u#h�kh�Yj jLh�kj�)`������u̃}� u-�j����    j jLh�kh lh�k�Ǟ����3��   �}�v�7����    3��~�} u�E   �URj ���P��E��MQ�URj���P��E��}� u:�}� @  w�M;M�w�u   ��t�U�U���� P�s�������败���0�E�^��]��������������������������������������������������������������������������U����E�����j j�E�Pj ���Q���t�}�u	�E�   ��E�    �E���]����������������������������U����E�E��M�Q�UR�EP�MQ�UR�EP�MQ�u^�����E��E�    �E���]��������������������������������U��E P�MQ�UR�EP�MQ�UR�EP������]������������������������U��j�h8�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t�}t	�E�    ��E�   �E܉E؃}� u#h��h�Yj jth�j�]������u̃}� u.�ԣ���    j jth�hTlh���1���������  �} t	�E�   ��E�    �UԉUЃ}� u#h��h�Yj juh�j�]������u̃}� u.�[����    j juh�hTlh��踛��������  j��]�����E�    �4��M��	�U�B�E�}� t�M�Q;Uu���}��   �}� tk�E�H���M̋U�ẺB�M̉M��}� uH�U�z t�E�H�U���M�9 t�U��M�Q�P��E�H�4�j�U�R��j�����<3�u&hزh�Yj h�   h�j�\������u��E������G����    ��   �}� tu�U�B���EȋM�UȉQ�EȉE��M�;4�tM�U�z t�E�H�U���M��E�H�J�U��    �E�4��H�4��E��M�4��h�   hD�jj�{W�����E�}� u�E�����薡���    �L�U��    �E�4��H�=4� t�4��E��M��A   �E�   �U�E�B�M�4��E������   �j�0�����ËE��M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��X!  迦�����3ŉE�ǅ����    ǅ����    ǅ����    �} u
�   �N  ������P�MQj�, ��u
ǅ����    �   i�  ������������  s��7���������Ƅ���� h  ������R������P���u8j h_  h�h�lh�lh4mh  ������Q薠����P��c����������������������P��������@vl������Q�������������D�������j hh  h�h�lh`�j�x�Q������������+й  +�Q������R�}d����P�Hc�����} t*�EP蔂������@v�MQ胂�����U�DÉ�����蓞���������膞���     �}uǅ����p��
ǅ�������   k� �M���t�E�������
ǅ�����Q�   k� �E���t�}uǅ�������
ǅ�������   k� �M���tǅ�������
ǅ�������} t�E�������
ǅ�����Q�} tǅ�������
ǅ�������} t�M�������
ǅ�����Q�} tǅ�������
ǅ������������ t�������������'�} t�E�������
ǅ�����Q������������������ tǅ����|��
ǅ�������} tǅ����Զ�
ǅ������������R������P������Q������R������P������Q������R������P������Q������R������P������Q�U��@lPhPmh�  h   ������Q�y����D������������ }*j h  h�h�lh��j"j�R����R�kS���� �B���������������� }8j h�  h�h�lh�h��h   ������R�ܜ����P�y`����h  h �������P�(u����������������uj�{c����j�sW��������u�   �3��M�3��t����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��|�]�������U��� ]������U���D ]������U��j�hX�h�Ld�    P���SVW���1E�3�P�E�d�    �E�E�}� ��  �M�y$ tj�U�B$P�6b�����M�y, tj�U�B,P�b�����M�y4 tj�U�B4P�b�����M�y< tj�U�B<P��a�����M�y@ tj�U�B@P��a�����M�yD tj�U�BDP�a�����M�yH tj�U�BHP�a�����M�y\�ytj�U�B\P�}a����j��S�����E�    �M�Qh�U܃}� t$�E܃����Iu�}�X�tj�U�R�9a�����E������   �j�؋�����j�jS�����E�   �E�Hl�M��}� t4�U�R�kg�����E�;4�t�}�8�t�M��9 u�U�R�xs�����E������   �j�k������j�E�P�`�����M�d�    Y_^[��]� ���������������������������������������������������������������������������������������������������������������������������������U��=|��t1�} u�|�P�Ej�����Ej �|�Q�6[�����UR�Շ��]������������������U��Q�s����E��}� u
j�e�����E���]��������������U����� �E��|�P��i�����E��}� uwj h  h,njh�  j�y�����E��}� tQ�M�Q�|�R�Z������t%j �E�P��f�����D �M���U��B�����j�E�P��^�����E�    �M�Q�X �E���]���������������������������������������������������U��j�h��h�Ld�    P��SVW���1E�3�P�E�d�    �E�@\�y�M�A    �U�B   �E�@p   �   k� �C   �Mf���   �   k� �C   �Uf���  �E�@hX��Mǁ�      j�[P�����E�    �U�Bh�   ���E������   �j萈�����j�"P�����E�   �U�E�Bl�M�yl u�U�4��Bl�M�QlR��b�����E������   �j�:�����ËM�d�    Y_^[��]���������������������������������������������������������������������������������U��Q�A����.�����u�Á��3��   h2\�H_�����|��=|��u	蜁��3��ijrh,njh�  j�f�����E��}� t�E�P�|�Q�X������u	�[���3��(j �U�R�Fd�����D �M���U��B�����   ��]��������������������������������������������������U��=|��t�|�P�{�����|������Ol��]����������������������U�졸�P� ]����������������U��} t#h`nh�Yj jWhxnj�M������u�j �&l����]�������������������������U��Qj��M�������P� �E��MQ� ���j�������E���]��������������������U��Q���P� �E��}� t�MQ�U�����u3���   ��]�����������������������������U��E���]����U��Q�E�����j j ���P�0 ��u�E������E���]��������������������U���*u��]�������U��Q�=�� u���j��u����h�   �u�����} t�E�E���E�   �M�Qj ���R�$��]����������������������������U��Q�E�    �}�wC�EP�i�����E��}� t�*�=�� u蛑���    ��MQ軃������u����UR襃�����l����    3���}� u�W����    �E���]������������������������������������������U��=�� u#h�rh�Yj jXh�rj�J������u̡��]���������������������������U���(����=�� u3���   ]���������������U�����    ]������������������U���SQ�E���E��EU�u�M�m���U��VW��_^��]�MU���   u�   Q�U��]Y[�� ��������������������U��j�h؈h�Ld�    P���SVW���1E�3�P�E�d�    �e���P� �E�}� t#�E�    �U��E�������   Ëe��E������-K���M�d�    Y_^[��]�����������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �e��4{���@x�E�}� t#�E�    �U��E�������   Ëe��E������g���M�d�    Y_^[��]�����������������������������������U��Q��z���@|�E��}� t�U��0J����]����������������U��h]'� ���]������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�x �Q  h (  h:^hJj �M��	Qj �o{�����E��}� u3��%  �U�R��q�����E�E�EԋM���M�}� v�U�U���� u�M�M�� ��j�nH�����E�    �U�z ��   j��k�����E܃}� ��   �E��P�k�����E؋M�U؉Q�}� t[j h�   hxsh�sht�E�P�M��Q�U�BP舎����P��Q�����M܋U�B��M܋U�B�A�M�U܉Q��E�P�t�����M�Q�h�����E������   �j������ËU�B�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������U��j�h8�h�Ld�    P���SVW���1E�3�P�E�d�    �E�x �f  j��F�����E�    �M�y �/  h (  j �U��	Rj 菏�����E��}� u"�E�    j��E�Ph��賓�����E��  �M�Q�o�����E�U�UЋE���E�}� v�M�M���� u�E�E��  ��j�i�����E܃}� ��   �E�    �M��Q�i�����E؃}� taj h  hxsh�thu�U�R�E��P�M�Q�l�����P�O�����U�E؉B�M܋U�B��M܋U�B�A�M�U܉Q��E�P�O}�����M�Q�C}�����E������   �j��}����ËU�B�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    j�D�����E�    �E�x ��   ����M��E�����U��U�}� t[�E�M�;Qu�E��M�Q�P�E�P�|�����4�M�M��U�z u#hDsh�Yj j9hxsj�0C������u�뙋M�QR��{�����E�@    �E������   �j�O|����ËM�d�    Y_^[��]����������������������������������������������������������������������U��j�hX�h�Ld�    P���SVW���1E�3�P�E�d�    j�ZC�����E�    �E�x ��   ����M��E�����U��U�}� t^�E�M�;Qu�E��M�Q�P�E�P�z�����7�M�M��U�z u&hDsh�Yj h�   hxsj��A������u�떋M�QR�tz�����E�@    �E������   �j��z����ËM�d�    Y_^[��]�����������������������������������������������������������������������������������U��j�hx�h�Ld�    P���SVW���1E�3�P�E�d�    j��A�����E�    �E�H�M��E�    ��U��U�}� t%�E�H�M��U�P�wy�����M�Q�ky�������E������   �j��y����ËM�d�    Y_^[��]��������������������������������������������������U���E��u	� (  f�M�URh:^hJ�EP�MQ�UR��s����]������������������������U��EP�MQ������]������������U��j �EP�MQ�UR�EP�MQ�UR��]����]����������U��Q�E�    �}et�}Eu%�E P�MQ�UR�EP�MQ�UR�:�����E��{�}fu!�E P�MQ�UR�EP�MQ脅�����E��T�}at�}Au%�U R�EP�MQ�UR�EP�MQ�:�����E��#�U R�EP�MQ�UR�EP�MQ�������E��E���]���������������������������������������������������U��j �EP�MQ�UR�EP�MQ�9����]��������������U���   �E�E��E��  �E�    �E�    �E�    �0   f�M��E�    �E�    3�f�U��E�    �E�    �E�    �E�    �EP��X�����G���} }�E    �} t	�E�   ��E�    �M��M��}� u&h�uh�Yj h�  h�uj��=������u̃}� uI�����    j h�  h�uh�wh�u�x|����ǅh���   ��X����W����h����L  �} v	�E�   ��E�    �E��E��}� u&hvh�Yj h�  h�uj�F=������u̃}� uC臃���    j h�  h�uh�whv��{�����E�   ��X����W���E��  �   k� �M� �U��9Uv	�E�   ��E�    �E��E��}� u&h�wh�Yj h�  h�uj�<������u̃}� uI����� "   j h�  h�uh�wh�w�<{����ǅt���"   ��X����gV����t����  �U܋�R�4��U��%�  �� �E��U��}��  �  �}� �  �}�u�E�E��	�M���M�j �UR�E�P�M��Q�UR�@D�����Eȃ}� t(�   k� �U�
 �EȉE���X�����U���E��w  �   ��U�
��-u�M�-�U���U�E� 0�M���M�} t�E�X��E�x�U�E��M���Mje�UR�[e�����E��}� t'�} t�E�P��E�p�E��M��U����U��E��  �MȉM���X����"U���E���  �U܋�R�?�T������ �E��U��E�E�t�M�-�U���U�E� 0�M���M�} t�E�X��E�x�U�E��M���M�} t�E�A��E�a�U��:�UċM܋�Q�4�&T��%�  �� �E��U��U�U�u[�E� 0�M���M�U܋�J���� ��x�����|�����x����|���u�E�    �E�    ��Ẽ��MЃ� �ẺM���U�1�E���E�M�M��U���U�} u�E��  ���X�����������   ��M����E܋�P���� ��l�����p�����p��� w��l��� �p  �E�   �E�    �M�EԋU��3����EԉU��E����   �} ~}�M܋�Q���� #E�#U��M���R��f�E��U���0f�U��E���9~�M�M�f�M��U�E���M���M�EԋUر�R���EԉU��U��f�U�E���E�q����M����   �U܋�R���� #E�#U��M��bR��f�E��E�����   �M�M��U����U��E����ft�U����Fu�M��0�U����U��ًE�;E�t/�M����9u�E���UčD�M����U�����M����U����U��E�����U��
�	�E���E�} ~�M�0�U���U���E����u�U��U�} t�E�P��E�p�E�M��U���U�M܋�Q�4�kQ��%�  �� +E�UЉE��U�}� |�}� r�U�+�E���E�"�M�-�U���U�E��؋M�� �ىE��M�U�U��E�� 0�}� |M	�}��  rBj h�  �M�Q�U�R�ل������0�M��U���Uj h�  �E�P�M�Q艄���E��U�U;U�u�}� |D�}�dr<j jd�E�P�M�Q脄���Ѓ�0�E��M���Mj jd�U�R�E�P�7����E��U�M;M�u�}� |D�}�
r<j j
�U�R�E�P�2����ȃ�0�U�
�E���Ej j
�M�Q�U�R�����E��U��E���0�M��U���U�E�  �E�    ��X����OP���E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�EP�MQ�!/����]��������������U���\�E�    �E P�M��=���} t	�E�   ��E�    �M��M�}� u&h�uh�Yj h�   h�uj�3������u̃}� u@��y���    j h�   h�uhvh�u�/r�����E�   �M��`M���E��\  �} v	�E�   ��E�    �E�E�}� u&hvh�Yj h�   h�uj�3������u̃}� u@�Gy���    j h�   h�uhvhv�q�����E�   �M���L���E���  �} ~�U�U���E�    �E���	9Ev	�E�   ��E�    �M܉M؃}� u&hHvh�Yj h  h�uj�^2������u̃}� u@�x��� "   j h  h�uhvhHv��p�����E�"   �M��*L���E��&  �E��tG�M�9-u	�E�   ��E�    �UUԉU��} ~	�E�   ��E�    �E�P�M�Q�w  ���U�U��E�8-u�M��-�U����U��} ~-�E��M��Q��E����E��M��~������   ��M����E��t	�E�    ��E�   �M�MM̉M��}�u�U�U���E�+E�M+ȉM�j h%  h�uhvh�vh�w�U�R�E�P�x����P��;�����M����M�} t�U��E�E����E��M�Q���0��   �M�Q���U�y�E��؉E��M��-�U����U��}�d|)�E���d   ���ЋE��ʋU��
�E���d   ���U��U����U��}�
|)�E���
   ���ЋE��ʋU��
�E���
   ���U��U����U��E��M��ЋE��� ���t �U����0uj�M��Q�U�R�8�����E�    �M���I���E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���\���3ŉE��E�E��M��M��E�    j�U�R�E�P�M��QR�P��A�����} t	�E�   ��E�    �M��M��}� u&h�uh�Yj hn  h�uj�^.������u̃}� u3�t���    j hn  h�uh�wh�u��l�����   �]  �} v	�E�   ��E�    �E��Ẽ}� u&hvh�Yj ho  h�uj��-������u̃}� u3�t���    j ho  h�uh�whv�xl�����   ��   �}�u�U�U��:�E܃8-u	�E�   ��E�    �} ~	�E�   ��E�    �M+M�+MĉMԋU܃:-u	�E�   ��E�    �} ~	�E�   ��E�    �E�P�M��Q�U�R�EE�E�P�J�����E��}� t�   k� �E� �E��(�MQj �U�R�EP�MQ�UR�EP��������E��E��M�3��K����]������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�EP�%r����]������������������U���@�E�H���M��UR�M��5���} t	�E�   ��E�    �E�E��}� u&h�uh�Yj h�  h�uj�+������u̃}� u@��q���    j h�  h�uhLxh�u�*j�����E�   �M��[E���E���  �} v	�E�   ��E�    �U�U�}� u&hvh�Yj h�  h�uj�+������u̃}� u@�Bq���    j h�  h�uhLxhv�i�����E�   �M���D���E��R  �M��tG�U�:-u	�E�   ��E�    �EE�E��M�;Mu�U�U��U��E�� 0�M����M��U�� �E�E��M�9-u�U��-�E����E��M�y j�U�R��
  ���E�� 0�M����M���U�E�B�E��} ��   j�M�Q�
  ���M��	w������   ��U����M����M��U�z }]�E��t�M�Q�ډU�&�E�H��9M}�U�U���E�H�ىM܋U܉U�EP�M�Q�;
  ���URj0�E�P�P�����E�    �M��vC���EЋ�]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���T���3ŉE��E�E��M��M��E�    j�U�R�E�P�M��QR�P�;�����} t	�E�   ��E�    �M̉Mă}� u&h�uh�Yj h�  h�uj�.(������u̃}� u3�on���    j h�  h�uhdxh�u��f�����   �*  �} v	�E�   ��E�    �E��E؃}� u&hvh�Yj h�  h�uj�'������u̃}� u3��m���    j h�  h�uhdxhv�Hf�����   �   �}�u�U�U��!�E܃8-u	�E�   ��E�    �M+MȉMԋU܃:-u	�E�   ��E�    �E�P�M܋UQR�E�P�MM�Q�D�����E��}� t�   k� �M� �E��$�URj �E�P�MQ�UR�EP��������E��E��M�3��E����]�����������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�EP�MQ�m����]��������������U���d���3ŉE��E�    �E�E��E� �M��M�j�U�R�E�P�M��QR�P��8�����} t	�E�   ��E�    �MĉM��}� u&h�uh�Yj h-  h�uj�z%������u̃}� u3�k���    j h-  h�uh|xh�u�d�����   �  �} v	�E�   ��E�    �ẺE��}� u&hvh�Yj h.  h�uj��$������u̃}� u3�:k���    j h.  h�uh|xhv�c�����   �9  �U܋B���EԋM܃9-u	�E�   ��E�    �UU��U؃}�u�E�E��!�M܃9-u	�E�   ��E�    �U+U��UȋE�P�MQ�U�R�E�P�GA�����EЃ}� t�   k� �E� �E��   �M܋Q��9U�}�E���E� �E�E�M܋Q���Uԃ}��|�E�;E|&�MQj�U�R�EP�MQ�UR�EP��������I�G�M��t!�U���E��M؃��M؃}� t��U��B� �EPj�M�Q�UR�EP�MQ�������M�3��AB����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP��I����]��������������U���V�EP�M��b,���M���t*�E�0�M��o������   ��;�t�U���U�̋E��M��U���U�}� ��   �E���t!�U���et�M���Et�E���E�ՋM�M��U���U�E���0u�U���U��E�0�M��o������   ��;�u	�U���U�E���E�M�U����M��U�E����E��}� t�ӍM��;��^��]����������������������������������������������������������������������������U��j �EP�MQ�UR�Af����]����������������������U����} t$�EP�MQ�U�R�K�����E�M��U��P��EP�MQ�U�R�`U�����E�M����]���������������������������������U��j �EP�f5����]��������������U����EP�M��C*���M�R��\������et�E���E�M�R�rm������u�E�Q�\������xu	�U���U�E��M��M��4m������   ��U���M���M�U��E��M�U���E��E��M��U��E���E�}� uҍM���9����]��������������������������������������������������������������U��Q�E�������Az	�E�   ��E�    �E���]������������������������U��} t#�EP�jI������P�MQ�UUR�'����]�������������������U��j jh�xhyh8yh   h   j �/����P�)����]����������������������������U��Q�E�    �	�E����E��}�
s�M���0�R� �M���0��ԋ�]��������������������U�����h���E��}� u3���  �E��H\Q�UR�  ���E��}� u	�E�    �	�E��H�M�}� u3��  �}�u�U��B    �   �  �}�u����t  �E��H`�M�U��E�B`�M��y�2  �Hz�U��	�E����E��HzLz9M�}kU��E��H\�D    �ҋU��Bd�E�M��9�  �u�U��Bd�   �   �E��8�  �u�M��Ad�   �   �U��:�  �u�E��@d�   �   �M��9�  �u�U��Bd�   �q�E��8�  �u�M��Ad�   �Z�U��:�  �u�E��@d�   �C�M��9�  �u�U��Bd�   �,�E��8� �u�M��Ad�   ��U��:� �u
�E��@d�   �M��QdRj�U���E��M�Hd��U��B    �E��HQ�U���U��E�B`�����]�������������������������������������������������������������������������������������������������������������������������������������������U��}csm�u�EP�MQ��0������3�]�������������U��Q�E�E��M��;Ut�E����E�k@zM9M�s��k@zU9U�s
�E��;Mt3���E���]�������������������������������U��E��]����U����E�    �=l� u�:���   i�  �M��}�  s���Y���U�Ƃ�� h  h��j �h���l;�����=(� t�(����t�(��U���E����E�E�M�Q�U�Rj j �E�P��   ���}����?s�}��r����w�M��U���;E�s����dh�   hpzj�M��U���P�u�����E�}� u����8�M�Q�U�R�E��M��R�E�P�M�Q�w   ���U�������E����3���]�������������������������������������������������������������������������������������������U��� �E�     �M�   �U�U��} t�E�M��U���U�E�    �E����"u/�}� u	�E�   ��E�    �U�U��E���M��U����U��w�E����U�
�} t�E�M����E���E�M���U��E����E��M�Q��&������t/�U����M��} t�U�E���
�U���U�E����E��M���t �}� �=����U��� t�E���	�'����M���u�U����U���} t�E�@� �E�    �M����t!�E���� t�U����	u�M����M��ߋU����u��  �} t�M�U��E���E�M����E��E�   �E�    �M����\u�E����E��M���M���U����"u`�E�3ҹ   ���uH�}� t�   �� �E����"u�U����U��#�E�    �}� u	�E�   ��E�    �E�E��M���M�U�U��E���E�}� t$�} t�M�\�U���U�E����U�
�ǋE����t�}� u�U���� t�M����	u�   �}� ��   �} tQ�E��Q��$������t)�U�E���
�U���U�E����E��M����E��M�U����M���M�)�U��P�$������t�M����M��U����M��U����M��U����U��_����} t�E�  �M���M�U����M�������} t�U�    �E���E�M����E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����=l� u�4���E�    ����E��}� u����e  �M����t,�E����=t	�U���U�E�P�?�����M��T�U���juh�zjj�E��P�2-�����E��M�� ��= � u�����   ����U��	�E�E��E��M������   �E�P�>�������E��M����=��   j~h�zjj�E�P�,�����M���U��: uj� �P��"����� �    ����rj h�   h�zh@{hX{�M�Q�U�R�E��Q�z[����P������U����U��B���j���P�i"�������    �M��    �p�   3���]�������������������������������������������������������������������������������������������������������U����E�    �E�    �=��N�@�t���%  ��t����щ���   �U�R�4�E�E��M�3M��M��D 3E��E��03E��E��U�R�,�E�3E�E��M�3M��M��U��E�3ЉU��}�N�@�u	�E�O�@���M���  ��u�U���G  ��U��U��E�����M��щ����]��������������������������������������������������������������������U����E�    �8�E��}� u3���   �E��E��M����t�E����E��M����u	�E����E��؋M�+M������M�j j j j �U�R�E�Pj j � �E��}� tjJh�{j�M�Q������E�}� u�U�R�<3��Dj j �E�P�M�Q�U�R�E�Pj j � ��uj�M�Q�������E�    �U�R�<�E��]���������������������������������������������������������������������������V�2��=�4s����t�Ѓ����4r�^������������V��5��=8s����t�Ѓ���8r�^������������U��EPj �MQ�UR�EP�R����]������������������U���@�E�    3��EĉEȉẺEЉEԉE؉E܍M��M��} t	�E�   ��E�    �U��U�}� u#h��h�Yj jph�{j��������u̃}� u.�'V���    j jph�{h,|h���N��������.  �} t�} u	�E�    ��E�   �M��M�}� u#hP|h�Yj jsh�{j�g������u̃}� u.�U���    j jsh�{h,|hP|�N��������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R��F�����E�} u�E��P�E��H���M�U��E�B�}� |!�M��� 3�%�   �E��M�����E����M�Qj ��M�����E��E��]���������������������������������������������������������������������������������������������������������������������������̀zuf��\���������?�f�?f��^���٭^�����|�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����|�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�����|���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-�|��p��� ƅp���
��
�t�������������������������������������������������������������������������������������������������������������������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�D>�����E�f�}t�m���������������������������������������������������ËT$��   ��f�T$�l$é   t�   ���|�   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �d��Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t���Z��=��Z��,$Z��}������������|�����   s��}��}������������|�����   v��}�����������������������������������������������������������������������������������������������������U��Q�E�   �} u�E�    �E���]������������������U��Q�E�   �} u�E�    �E���]������������������U��Q�E�   �} u�E�    �E���]������������������U��3�]����������U��j�h8�h�Ld�    P��SVW���1E�3�P�E�d�    �=4�8�tAj�n	�����E�    h8�h4���J�����4��E������   �j�A����ËM�d�    Y_^[��]��������������������������������������������������U�� �]�������U���]�������U����} u3��   jU�EP�D�����E��}�Ur3��ihw  h�j�M��T	R������E��}� u3��@j hz  h0h̑h ��E���P�MQ�U���R�E�P�����P������E���]������������������������������������������������������U��EP�MQ� =����]������������U��EP�*����]����������������U������]�������U��j hc  h0h �h@��EP�MQ�UR�M����P�[�����   k� �U��
�   ��t!�M���   Qhđj�UR�EP��+�����   k� �E��   ��t!�U��   Rhȑj�EP�MQ�+����]���������������������������������������������������������U���h�  j �EP��,�����M���u3���  �   k� �U�
��.up�   �� �U�
��t]j h9  h0h�h0�j�   �� MQj�U��   R�����P������   k�3ҋEf��   3��j  �E�    �	�M���M�h4��UR��L�����E��}� u����6  �E��Mf�Af�U��}� uI�}�@sC�E���.t:j hG  h0h�h@��M�Q�URj@�EP�`����P�w�����   �}�uL�}�@sF�M���_t=j hJ  h0h�h8��U�R�EPj@�M���   Q�����P�"�����^�}�uS�}�sM�U���t	�E���,u<j hM  h0h�h(��M�Q�URj�E   P�����P�����������)�M���,u��U���u��E��M�TA�U����3���]�����������������������������������������������������������������������������������������������������������������������������������������������������U����q5���E��E��Hp��u	�E�   ��E�   �U�U�E�E��M����M��}�wC�U��$�h#�E��Hp���U��Jp�   �E��Hp����U��Jp�   �   � ������z3�t	�E�   ��E�    �M��M�}� u&h�~h�Yj h�   h0j�h������u̃}� u.�H���    j h�   h0h�h�~�A���������E��]��"�"�"�"������������������������������������������������������������������������U��VW�} t0�} t*�E;Et"�.   �u�}�M�    �UR�����_^]������������������U���  ���3ŉE��} |�}�} u3��7h�   ������Pj��MQj j � ��u3��������R�EP�5�����M�3�������]�����������������������������������U���  ���3ŉE��$3���   ��(�����(������� �����(����������ǅ����   ��(�����"  ��$���ǅ����   ǅ,���    ǅ���    �} u3��T  j h�  h0hT�hx�jU��(���P  P�MQ�UR������P��
�����E���Cu^�   �� �E���uKj h�  h0hT�h�hp��UR�EP�G����P�
�����} t	�M�    �E�  �UR�m)������,�����,����   s6�EP��$���Q�*�������  �UR�����P��)�������  ǅ������ǅ ���    ǅ���    ǅ���   �   k�����3�������t
ǅ���    �MQ��0���R��7������uQ����� t%��0���P�� ���Q��0���R��)����������#��0���P�� ���Q��0���R�R(�������������� tq��0���P�����Q��$���R��M�����} tIj h�  h0hT�hx���P���P�(������P��P���Q�UR�EP������P�	�����m  �MQ��G�������  j�����Rh  �EP� �������t	����� u������������� ����
j h�  h0hT�hp���,�����P�MQ�����R��$���P�_����P�v����j h�  h0hT�h���,�����Q�UR�EP�MQ�"����P�9����j h�  h0hT�h����,�����R�EPjU��(�����P  Q������P�������Qj h  h0hT�hp��UR�&������P�EPjU��(�����P  Q�����P�����3��   �U���tQ��,����   sEj h  h0hT�h ���,�����Q�UR�����P�����Q�2����P�I�����3ҋ����f��} tj�� ���Q�UR�����j h  h0hT�h����$���P�MQ�UR�NC����P��������$����M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hȉh�Ld�    P��SVW���1E�3�P�E�d�    �} ��   j�p������E�    �E�x t-�M�Q�����Hu�M�yX�tj�U�BP�������E������   �j�~3����ËM�9 tcj�������E�   �U�P������M�9 t#�U��8 u�M�98�t�U�P� �����E������   �j�3�����j�MQ�M�����M�d�    Y_^[��]����������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �`+���E�h�  h�jjj�l�����E�}� u�<?���    3��   ��3���7���E�M��Ql��E�M��Qh�Pj�������E�    �E�Q������E������   �j��1�����j�o������E�   �U�B�   ���E������   �j�1����ËE�M�d�    Y_^[��]������������������������������������������������������������������������U����E�    �} |�}�} u3��  hL  h�jjj�%�����E��}� u��=���    3��  hQ  h�jjh�   �������E��E��M���}� u j�U�R�������=���    3��=  hW  h�jjh   ������E�E��M�H�}� u0j�U��P�����j�M�Q������L=���    3���   h8��U��P�������MQ�UR�E��Q�x	  ����uDj�U��BP�P�����M��R������E��Q������j�U�R�&�����E�    �l�E��HQ�U���HQ��������tDj�U��BP�������M��R�Y�����E��Q�����j�U�R�������E�    ��E��H�   �E���]���������������������������������������������������������������������������������������������������������������������������U����E�E��E�    �	�M����M��U�;U}A�E����E�j h&  h0h �h8��M��Q�R�EP�MQ�6=����P���������E�    ��]�������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} |�}	�E�   ��E�    �E؉Eԃ}� u&h�h�Yj h  h0j�y�������u̃}� u0�:���    j h  h0h`�h��3����3��  �&���E��$/���U��Bp���M��Ap�E�    h  h�jjh�   �s�����E�}� �  j��������E�   �U��BlP�M�Q�������E�    �   �j�-����Ã}� ��   �UR�EP�M�Q�K  ���E܃}� ��   �} th���UR��������t
��   j�P������E�   �E�P�M���lQ��5�����U�R�M�����E��Hp��u$� ���u�E��HlQh4��5�����g  �E�    �   �j�F,�������U�R�������E�P� �����E������   ��M��Qp���E��PpËE܋M�d�    Y_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�   �E�    �E�    �E�    �E�    �E�  hd  h�j�E�P��������E�}� u3��X  �M���M��U�����U�3��M�f��U��   �E�   �	�E����E��M����U�D
Ph�kM���8}Rj�E�P�M�Q�������}�}kj hp  h0h�h�h���U�R�E�P�9����P��������M������U�D
P�M����U�D
P�U������t�E�    �{  �}� �/  �   k� �E�| tZ�   k� �E�L�����JuA3�u#j h�Yj hy  h0j�y�������u�j�   k� �M�TR��������   k� �U�|
 tZ�   k� �U�D
�����IuA3�u#j h�Yj h~  h0j��������u�j�   k� �E�LQ�������   k� �M�D    �   k� �M�D    �   k� �M�U�T�   k� �U�E��D
�E��L  �B  j�M�Q�)������   k� �M�| tZ�   k� �M�T�����HuA3�u#j h�Yj h�  h0j�<�������u�j�   k� �U�D
P�������   k� �E�| tZ�   k� �E�L�����JuA3�u#j h�Yj h�  h0j���������u�j�   k� �M�TR�Q������   k� �U�D
    �   k� �U�D
    �   k� �U�D
    �   k� �U�D
    �   ���M�D��������]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����  ���3ŉE��} tF�} t�EP�MQ�UR�0  ����,�����E���M�T��,�����,�����0�����  ǅ ���   ǅ4���    �} ��  �   k� �E���L�a  �   �� �E���C�I  �   ��E���_�2  �U��<���h|���<���P�s(������@�����@��� t$��@���+�<�������8���t��@������;u3��  ǅD���   ���D�������D�����D���J��8���R��<���Pk�D�����8}R�I4������u k�D�����8}Q�����9�8���u�랋�@�������@���h����@���P�3������8�����8��� u��@������;t3��f  ��D�����   j h�  h0h��h����8���P��@���Qh�   ������R������P��������8�������$�����$���  s���)��3ɋ�$���f������������P��D���Q�UR��  ����t��4�������4�����8�����@����J��<�����<������t��<�������<�����<������������4��� t�EP������������
ǅ���    �������0����&  j jU��H���Rh�   ������P�MQ��+������0�����0��� ��   ǅD���    ���D�������D�����D���|��D��� tn��D������M�TR������P�L������t;������Q��D���R�EP��  ����t��4�������4����
ǅ ���    ���4�������4����l����� ��� t�EP�r�������0����3��4��� t�MQ�U�������(����
ǅ(���    ��(�����0�����EP�)�������0�����0����M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����  ���3ŉE�Vǅ<���    ǅ4���    ǅ$���    ��������������  ��D���ǅ(���   �� ���QjU��H���Rh�   ������P�MQ� )������u3��<  �U���E�LQ������R�������u�E���M�D�	  ������R����������$���h�  h�j��$����L Q��������<�����<��� u3��  ��<�������4����E���M�T������E�M����   ������E�H�����j h�  h0hT�h��������R��$���P��4���Q�-����P�9������U���E��4����L�   k� ��������Cu'�   �� ��������u�M�UǄ��       ���H���P������M�U����   �}�:  �E�� ����H��(�����D����L���T����,�����0���ǅ@���    ���@�������@�����@���;�(�����   �U��@�����D����R;�uT��@��� tG��@�����D������D��   k� ��D�����D��@�����D�����,����Ћ�0����L��]�V��@�����D����ЋT�������������@�����D�����,�������0����T��������,����������0���������@���;�(�����   j�E�HQ������Rjh ~jj �p��������   ǅ8���    ���8�������8�����8���s$��8�����M�������  ��8���f��E������h�   �`�Q������R�W�������u�   k� ��D����D
   ��   k� ��D����D
    ��   k� ��D����D
    �   k� ��D����E�@�
�   k� �E��D����T�Pp�&�}u�E�� ����H��}u�U�� ����B�MQkU��@}�Ѓ���tb�M���U������D
j�M�U����   P��������M�U���������   j��<���Q��������U������B3���   ���������   �M���U�D
�����I��   3�u#j h�Yj hH  h0j���������u�j�M���U�D
P�P�����j�M���U�D
P�8�����j�M�U����   P� ������M���U�D
    �E�MǄ��       ��<��� t��<����   �E���M��<����T�E���M�D^�M�3��� ����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��4����   � ��4����   ���4��Qt���]���������������������������U����E�    �} u�E��Q�U�}  t	�E�	   ��E�   j j �EP�MQ�U�R�EP� �E��}� u3���   3�uS�}� ~M�}����wD�U���R�2�������t#h��  �E��L Q��	����P�{!�����E���E�    �U��U���E�    �E�E��}� u3��a�M���Qj �U�R������E�P�M�Q�UR�EPj�MQ� �E�}� t�UR�E�P�M�Q�UR� �E�E�P��������E��]��������������������������������������������������������������������������������U����EP�M������M Q�UR�EP�MQ�UR�EP�M��+��P�H������E��M������E���]��������������������U��EP�MQ�UR�EP�����]��������������������U���T�E�    �} t�} u3��`  �} t�} v3��Mf��} t	�E�   ��E�    �U��U�}� u#h|�h�Yj jEh��j���������u̃}� u.�$���    j jEh��h�h|��j���������  �MQ�M��L����} �  �M��*����   �����    uj�M�;MsG�UU�f��Mf��UU����u�M��M�M��>����E��g  �U����U��E���E뱋M��M�M������E��=  �  �UR�EPj��MQj	�M���)����BP� �E��}� t�M����M��M�������E���  �� ��zt*��"��� *   3ҋEf��E������M������E��  �M�M�U�U��	�E����E��M�M؋U���U�}� ts�E����ti�M��R)��P�U��P�b*������tH�   �� �U��
��u,�d"��� *   3ɋUf�
�E������M������E��.  �	�E����E��o����M�+M�MЋUR�EP�M�Q�URj�M���(��� �HQ� �E��}� u*��!��� *   3ҋEf��E������M������E��   �M��MȍM��}����E��   �   �M��l(����   �����    u�MQ�i�����EčM��>����E��j�`j j j��URj	�M��'(��� �HQ� �E��}� u!�K!��� *   �E������M�������E�� ��U����U��M�������E���M��������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���T�E�    �} u�} t�} t�} w	�E�    ��E�   �E��E�}� u&h8�h�Yj h�   h��j�n�������u̃}� u3����    j h�   h��h�h8��	�����   �  �} tY3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E��M���Qh�   �U��R��������} t	�E�     �MQ�M��{����U;Uv�E�E���M�M�U�U��}����w	�E�   ��E�    �E�E�}� u&h�h�Yj h  h��j�T�������u̃}� u@����    j h  h��h�h��������E�   �M�� ����E���  �M��%��P�U�R�EP�MQ������E��}��uy�} tY3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E܋M���Qh�   �U��R����������� �EčM������E��G  �M����M��} �  �U�;U��   �}���   3��Mf��}�tJ�}���tA�}v;�U��9h�s
�h��E��	�M���M؋U���Rh�   �E��P��������M�;Mw	�E�   ��E�    �UԉUЃ}� u&h<�h�Yj h  h��j��������u̃}� u=����� "   j h  h��h�h<��?�����E�"   �M��p����E��9�M�M��E�P   3ҋE��Mf�TA��} t�U�E���M̉M��M��5����E���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��=� uh��EP�MQ�UR�K�������j �EP�MQ�UR�1�����]��������������������������������U��j �EP�MQ�UR�EP�MQ������]��������������U����E���E��M�M��U����U�t�E����t�U����U����}� t�E����u�E�+E������E��]������������������������U��EP�MQ�UR�EP�������]��������������������U���   ���3ŉE��E�    �E�    �} t�} u3���  �} t	�E�   ��E�    �EĉEȃ}� u#ht�h�Yj jfh��j��������u̃}� u.�����    j jfh��h�ht��*��������M  �UR�M������} �9  �M��H ��� �   �ჼ�    ��   �U�;Usv�E����   ~"�T��� *   �E������M�������E���  �UU��E��
�U��E��M���M�}� u�U��U��M�������E��  �E����E�낋M��M��M������E��  �|  �M������zt��   �} v�EP�MQ�������E�U�Rj �EP�MQ�UR�EPj �M��K����QR� �E��}� t3�}� u-�EE��H���u	�U����U��E��E��M������E���  �<��� *   �E������M�������E���  ��  �M�Qj �UR�EPj��MQj �M������BP� �E��}� t�}� u�M����M��M������E��q  �}� u�� ��zt"���� *   �E������M��[����E��>  �U�;U�  �E�Pj �M��=����QtR�E�Pj�MQj �M��#����BP� �E؃}� t�}� t"�A��� *   �E������M�������E���  �}� |�}�v"���� *   �E������M������E��  �M�M�;Mv�U��U��M������E��~  �E�    ��EЃ��EЋM����M��U�;U�}4�EE��MЊT��EE����u�U��U��M��F����E��)  벋E���E������M��M��M�� ����E��  ��   �M������   �����    uq�E�    �M�M��	�Uԃ��UԋE����t:�U��=�   ~"���� *   �E������M������E��   �M̃��M�볋ỦU��M������E��t�j�E�Pj j j j��MQj �M��q����BP� �E��}� t�}� t���� *   �E������M��8����E���M����M��M��"����E���M������M�3��������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���4�E�    �} t�} w�} u�} t	�E�    ��E�   �E��E�}� u&h8�h�Yj h@  h��j�N�������u̃}� u3����    j h@  h��h��h8��������   �  �} tU�U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U��E�Ph�   �M��Q��������} t	�U�    �E;Ev�M�M���U�U�E�E��}����w	�E�   ��E�    �M�M�}� u&h�h�Yj hL  h��j�D�������u̃}� u3����    j hL  h��h��h���
�����   �  �EP�M�Q�UR�EP��������E��}��uf�} tT�M� �}�tH�}���t?�}v9�U��9h�s
�h��E��	�M���M܋U�Rh�   �E��P����������� �&  �M����M��} �  �U�;U��   �}���   �E�  �}�tI�}���t@�}v:�M��9h�s�h��U��	�E���E؋M�Qh�   �U��R�������E;E�v	�E�   ��E�    �MԉMЃ}� u&h�h�Yj hd  h��j��������u̃}� u0����� "   j hd  h��h��h��W	�����"   �(�E�E��E�P   �MM��A� �} t�U�E���E̋�]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�<�����]����������������������U��j �EP�MQ�UR�EP�MQ�f�����]��������������U��j�hX�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j��������E�    �E�    �	�E���E�M�;���N  �U�|��<� ��   �M�|����H��   ��   �U�|����Q�� �  ��   �}�~�}�}�E��P�������u��   �M�|���P�M�Q��������U�|����Q��   t�E�|���R�E�P�������0����M�|����E��   �{jZh8�jj8��������E܋M�|��E܉��}� tNj h�  �M�|����� P�������M�|����� P�  �M�|����E��M��A    ������}� tB�U��B% �  �M��A�U��B    �E��@    �M��    �U��B    �E��@�����E������   �j�P ����ËE��M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������������������������������������������������U���X�E�    ���E��E�    �E�    �E�    �} u#h��h�Yj jDh��j��������u̃} u#h�h�Yj jEh��j���������u̃} u#ht�h�Yj jFh��j��������u̋M��� u�E���E��M��U��}�at8�}�rt�}�wt�<�E�    �E����E��   �E�  �M����M��   �E�	  �U����U��v3�t	�E�   ��E�    �M܉M؃}� u#h8�h�Yj jbh��j���������u̃}� u-�@���    j jbh��h��h8������3���  �E�   �E���E�M����<  �}� �2  �E��M�U�� �U�}�T��  �E����f�$��f��  �U���t	�E�    �'�E����E��M�����M��U��ʀ   �U��E�����E��  �M��� �  t	�E�    ��U��� �  �U��  �E�% �  t	�E�    ��M��� @  �M��u  �}� t	�E�    ��E�   �U��� @  �U��N  �}� t	�E�    ��E�   �E�%�����E��(  �}� t	�E�    ��E�   �M��� �M��  �}� t	�E�    ��E�   �U����U���   �E�%   t	�E�    ��M���   �M��   �U���@t	�E�    �	�E���@�E��   �M��ɀ   �M��   �E�   �E�    �|3�t	�E�   ��E�    �EԉEЃ}� u&h8�h�Yj h�   h��j��������u̃}� u0�����    j h�   h��h��h8��H����3��  �����}� �w  �U��� u�M���M��j�URhh��/������t|3�t	�E�   ��E�    �MȉMă}� u&h8�h�Yj h�   h��j���������u̃}� u0�6���    j h�   h��h��h8�� ����3���  �E���E�M��� u�E���E��M���=t|3�t	�E�   ��E�    �M��M��}� u&h8�h�Yj h�   h��j�O�������u̃}� u0����    j h�   h��h��h8��������3��1  �E���E�M��� u�E���E��jhl��MQ�K�������u�U���U�E�   �E���   jht��MQ��������u�U���U�E�   �E��   jh���MQ���������u�U���U�E�   �E��|3�t	�E�   ��E�    �U��U��}� u&h8�h�Yj h  h��j�'�������u̃}� u0�h���    j h  h��h��h8��������3��	  �M��� u�E���E��M���u	�E�   ��E�    �E��E��}� u&h��h�Yj h  h��j菿������u̃}� u-�����    j h  h��h��h���*�����3��th�  �UR�E�P�MQ�U�R��������t3��O�\����\��M�M��U��E��B�M��A    �U��    �E��@    �M��A    �U��E��B�E���]ÍI a#a�bbb�bb�a>b`a�a�a�a�b 	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������SVW�T$�D$�L$URPQQh�id�5    ���3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�c����   �C�*����d�    ��_^[ËL$�A   �   t3�D$�H3��i���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�����3�3�3�3�3���U��SVWj RhvjQ�5���_^[]�U�l$RQ�t$������]� ����������������������������������������������������������������������������������������������U��H  �o�����3ŉE��} tǅ����   �
ǅ����    ������������������ u#h��h�Yj j\hȗj�:�������u̃����� u.�x ���    j j\hȗh8�h�������������  �U������������P�\������������������y }�������B    jj ������P������������������ }����  ��������������������0��L$�����������������B%  u������������+A�Y  �������������
+H�������������B����  ���������_  ��������������������0��|0 �8  �������������
+H�鉍�����������z u��������  �  j ��������������������0��D
,P�L
(Q������R��������������������������������������0�������������������������������;T(u������������������;T,t����!  j ������Ph   ������Q��������������������0��R�� ��u�����  j ������P������Q��������}����  ������;�����v����  �������������������������������������������� ��   ������������9�����ss���������u5������������9�����s�������H��
u������������������������X���������������������������P���������������+ʋ�3�������������  ��������������������0��T��   tO�������H���������������������������������;s���������
u�����������������#�������B%�   u�y����    ����$  ������ u�������  �������Q����  �������x uǅ����    �  �������������+B������A��������������������������0��T��   �^  jj ������P�p�����;�������   �������Q������������������H���������������������������;�����s���������
u���������������ċ������Q��    t���������������   j ������Q������R���������}�����   ������   w*�������H��t�������B%   uǅ����   ��������Q��������������������������0��D
��t����������������������u�������艅����������+�������������������u�������艅����������������M�3�������]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hx�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h �h�Yj j0hȗj蹱������u̃}� u+������    j j0hȗh(�h ��W���������@�UR��������E�    �EP��������E��E������   ��MQ�|�����ËE܋M�d�    Y_^[��]������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u������     ������ 	   �����  �} |�E;<�s	�E�   ��E�    �M��M܃}� u#hMh�Yj jAh`�j�J�������u̃}� u9膵���     ����� 	   j jAh`�h��hM�����������L  �E���M������0��D
��t	�E�   ��E�    �M؉Mԃ}� u#h�Mh�Yj jBh`�j謯������u̃}� u9�����     ������ 	   j jBh`�h��h�M�?���������   �EP�������E�    �M���U������0��L��t�UR�EP�MQ�������E��D�h���� 	   �X����     �E�����3�u#h(Nh�Yj jMh`�j�ݮ������u��E������   ��MQ般����ËE�M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������U����EP�ڷ�����E��}��u:�A���� 	   3�u#hИh�Yj jkh`�j�ȭ������u̃����   �E�    �E�    j�E�P�M�Q�U�R�E�P�� ��u�� P�U���������   �E��E�U��MQ�U�R�E�P�M�Q�U�R�� ��u�� P����������g�}� t&j j �E�P�M�Q�U�R�� �n����    ����;�E���M������0��D
����M���U������0��D�E��]������������������������������������������������������������������������������������U���X�E�    ���E��E�    �E�    �E�    �} u#h��h�Yj jDh��j�2�������u̃} u#h�h�Yj jEh��j�	�������u̃} u#ht�h�Yj jFh��j��������u̋M��� u�E���E��M��U��}�at8�}�rt�}�wt�<�E�    �E����E��   �E�  �M����M��   �E�	  �U����U��v3�t	�E�   ��E�    �M܉M؃}� u#h8�h�Yj jbh��j�.�������u̃}� u-�o����    j jbh��h\�h8��������3���  �E�   �E���E�M����<  �}� �2  �E��M�U�� �U�}�T��  �E������$�����  �U���t	�E�    �'�E����E��M�����M��U��ʀ   �U��E�����E��  �M��� �  t	�E�    ��U��� �  �U��  �E�% �  t	�E�    ��M��� @  �M��u  �}� t	�E�    ��E�   �U��� @  �U��N  �}� t	�E�    ��E�   �E�%�����E��(  �}� t	�E�    ��E�   �M��� �M��  �}� t	�E�    ��E�   �U����U���   �E�%   t	�E�    ��M���   �M��   �U���@t	�E�    �	�E���@�E��   �M��ɀ   �M��   �E�   �E�    �|3�t	�E�   ��E�    �EԉEЃ}� u&h8�h�Yj h�   h��j�ܨ������u̃}� u0�����    j h�   h��h\�h8��w�����3��  �����}� �w  �U��� u�M���M��j�URh����������t|3�t	�E�   ��E�    �MȉMă}� u&h8�h�Yj h�   h��j�$�������u̃}� u0�e����    j h�   h��h\�h8�������3���  �E���E�M��� u�E���E��M���=t|3�t	�E�   ��E�    �M��M��}� u&h8�h�Yj h�   h��j�~�������u̃}� u0�����    j h�   h��h\�h8�������3��1  �E���E�M��� u�E���E��jh ��MQ��������u�U��
�U�E�   �E���   jh,��MQ�X�������u�U���U�E�   �E��   jh@��MQ�(�������u�U���U�E�   �E��|3�t	�E�   ��E�    �U��U��}� u&h8�h�Yj h  h��j�V�������u̃}� u0�����    j h  h��h\�h8��������3��	  �M��� u�E���E��M���u	�E�   ��E�    �E��E��}� u&h��h�Yj h  h��j辥������u̃}� u-������    j h  h��h\�h���Y�����3��th�  �UR�E�P�MQ�U�R�O�������t3��O�\����\��M�M��U��E��B�M��A    �U��    �E��@    �M��A    �U��E��B�E���]Ë��z�zc|3|R|�{�{|1{z{�{V{s| 	
�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U������]��E�E��M������U�ҁ�   �ʉM��E���]����������������U������]��E�E��M��M�U��%����M���ҁ�   �M��E���]���������������������U������]��E�E��M������U��   �ʉM��E���]������������������U������]��E�E��M�M�U��U��E��������U�%   �ȋU��
�E���]�����������������U���E%�  =�  u3���   ]�������������������U����E%�  =�  uP���E�$��������E��}�t�}�t�}�t��   �   �   �   �   �   �   �   �M�� �  �M��U���  u+�E����u�} t�}� t	�E�   ��E�   �E��B�E��������Dz�}� t	�E�    ��E�@   �E���}� t	�E�   ��E�   �E��]�����������������������������������������������������������������U���E%�  =�  u�M����u�} u�U���  ���  u�   �3�]�����������������U������]�h��  h?  �������E��E%�  =�  ��   ���E�$�I������E��}� ~C�}�~�}�t�5h��  �M�Q�5������E�   �U�R���E�$j%�������   �E�P�E��`���$���E�$j%j�$������q�E��������Dz)�M�Q�p������$���E�$j%j�������:�U�R���E�$������؃��E���E��E��]�h��  �M�Q�y������E��]���������������������������������������������������������������������������������U���$���]�h��  h?  �������E��E%�  =�  t�M���  ���  ��   �U���  ���  u�E����u(�} u"�M���  ���  uC�U����u�} t3�E�P�E�E���$���E�$���E�$j&j蹜����$�\  �M���  ���  t�U���  ���  u%�E�P���E�$���E�$j&�������  �E�E������Dzh��  �M�Q��������E��  �E��������Dz$�E�   �E�]����z	�E�    ��E�   ����]����z�E�]����At���]����Au-�E�]����z �U���U�E�E��} u	�M����M��P���]����z�E�]����{���]����Au+�E�]����Au�U���U�E�E��}� u	�M����M��U���  uv�E�����u�}� tf�M�Q���E��$�J������]�U���   R���E��$�L������]�E�P���E��$���E�$���E�$j&j������$�   �}�  �u�}� t�}�  ��ui�}� uc�M�Q���E��$��������]܋U��   R���E��$�ȴ�����]�E�P���E��$���E�$���E�$j&j�n�����$�h��  �M�Q�������E��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EP���E�$�w�����]�������U��EPj �MQh�]�8�����]���������������������U���0�E�    3��EԉE؉E܉E��E�E�E�MЉM��} t	�E�   ��E�    �U��U�}� u&h��h�Yj h�  h�{j胙������u̃}� u.������    j h�  h�{h��h������������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]��������������������������������������������������������������������U��EP�MQ�URh�]�������]�������������������U��EPj �MQh_a������]���������������������U��EP�MQ�URh_a�v�����]�������������������U���@�E�    3��EĉEȉẺEЉEԉE؉E܍M��M��} t	�E�   ��E�    �U��U�}� u#h��h�Yj jph�{j�Ɨ������u̃}� u.�����    j jph�{hx�h���d���������  �} t	�E�   ��E�    �M��M�}� u#hX�h�Yj juh�{j�M�������u̃}� u.�����    j juh�{hx�hX������������   �E��@����M��AB   �U��E�B�M��U��EP�MQ�UR�E�P��������E�} u�E��Q�M��Q���U�E��M�H�}� |"�U���  3Ɂ��   �M��U�����M����U�Rj ��������E��E��]���������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR������]����������������������U����EPj �MQ�UR�EPh�]諷�����E��}� }	�E�������M��M��E���]�����������������������������U����EP�MQ�UR�EP�MQh�]�I������E��}� }	�E�������U��U��E���]���������������������������U���@�E�    3��EĉEȉẺEЉEԉE؉E܍M��M��} t	�E�   ��E�    �U�U��}� u#h��h�Yj jph�{j覔������u̃}� u.������    j jph�{h��h���D���������W  �} t�} u	�E�    ��E�   �M�M�}� u#hP|h�Yj jsh�{j�'�������u̃}� u.�h����    j jsh�{h��hP|������������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R�U���E��} u�E��{�}� |X�E��H���M�U��E�B�}� |!�M��� 3�%�   �E��M�����E����M�Qj �������E��}��t�E���UU�B� �E��x }�����������]�����������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP�MQ������]��������������U���0�E������E�    �} t	�E�   ��E�    �E�E��}� u&h�h�Yj h  h�{j�	�������u̃}� u1�J����    j h  h�{hȚh�����������'  �} u�} u�} u3��  �} t�} v	�E�   ��E�    �U�U�}� u&h8�h�Yj h  h�{j�k�������u̃}� u1�����    j h  h�{hȚh8�����������  �M;M��   �o�����U��EP�MQ�UR�E��P�MQhL`��������E��}��u~�}�t\�}���tS�U��;UsH�E���M+�9h�s�h��U���E���M+ȉM�U�Rh�   �E�M�TR螷����������8"u
������M�������  �`������U��EP�MQ�UR�EP�MQhL`�A������E��UU�B� �}��u"�}�u�t����8"u
�j����M������f  �}� ��   �   k� �M� �}�tH�}���t?�}v9�U��9h�s
�h��E��	�M���M��U�Rh�   �E��P蹶�����}��uz3�t	�E�   ��E�    �U܉U؃}� u&h��h�Yj hB  h�{j�^�������u̃}� u.����� "   j hB  h�{hȚh�����������������z�}�t\�}���tS�M���;MsH�U����E+�9h�s�h��M���U����E+EԋM�Qh�   �U��E�LQ�ҵ�����}� }	�E�������U��UЋEЋ�]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EPj �MQ�UR�EPh_a苯�����E��}� }	�E�������M��M��E���]�����������������������������U����EP�MQ�UR�EP�MQh_a�)������E��}� }	�E�������U��U��E���]���������������������������U���$�E������} t	�E�   ��E�    �E��E�}� u&h�h�Yj h�   h�{j蠌������u̃}� u1������    j h�   h�{h�h��;����������  �} t�} v	�E�   ��E�    �U��U�}� u&h8�h�Yj h�   h�{j��������u̃}� u1�\����    j h�   h�{h�h8�����������s  �MQ�UR�EP�MQ�URhL`辭�����E��}� }^�   k� �U�
 �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U�E�Ph�   �M��Q�k������}��uz3�t	�E�   ��E�    �E�E��}� u&h��h�Yj h�   h�{j��������u̃}� u.�Q���� "   j h�   h�{h�h������������k�}� |b�}�t\�}���tS�U���;UsH�E����M+�9h�s�h��U���E����M+ȉM܋U�Rh�   �E��M�TR胱�����E���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP������]������������������U���8  ���3ŉE�ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    �EP�� ����ْ��ǅ����    �V�����d����} tǅ���   �
ǅ���    �������$�����$��� u&h �h�Yj h  hx�j譈������u̃�$��� uI������    j h  hx�h؛h ��E�����ǅ���������� ����p����������W  �E��\�����\����Q��@��   ��\���P袻�����������������t-�������t$�������������������0�������
ǅ����������H$�����х�uV�������t-�������t$�������������������0���0����
ǅ0������0����B$�� ���ȅ�tǅ,���    �
ǅ,���   ��,�����P�����P��� u&hp�h�Yj h	  hx�j�0�������u̃�P��� uI�n����    j h	  hx�h؛hp��������ǅ���������� ���������������  �} tǅ���   �
ǅ���    �������H�����H��� u&h��h�Yj h  hx�j臆������u̃�H��� uI������    j h  hx�h؛h��������ǅ���������� ����J����������1  ǅ����    ǅ����    ǅ����    ǅ����    ǅ|���    �E��������������������E���E������ ��  ������ ��  �������� |%��������x�������������(����
ǅ(���    ��(�����������������������������������������@�����@����%  ��@����$���ǅ����    �� ����7���P������R�F���������   ������P�MQ������R�3  ���E��������U���U��������tǅ���   �
ǅ���    �������8�����8��� u&h�h�Yj h�  hx�j腄������u̃�8��� uI������    j h�  hx�h؛h�������ǅ���������� ����H����������/  ������P�MQ������R�V  ����  ǅ����    ������������������������������������ǅ����    ǅ��������ǅ����    �  �������������������� ������������wj��������ر�$������������������E���������������4���������������#�������ɀ   ����������������������  ��������*u:�MQ������������������ }���������������������؉������k�����
�������DЉ������  ǅ����    �  ��������*u'�UR�x����������������� }
ǅ���������k�����
�������TЉ������F  ��������������������I������������.�3  �������� ��$���M���lu�E���E��������   �����������������������   �E���6u,�U�B��4u �M���M�������� �  �������   �E���3u)�U�B��2u�M���M������������������S�E���dt7�U���it,�M���ot!�E���ut�U���xt�M���Xu�ǅ����    ������#�������� ���������������   ��������  ��������������������A������������7�)
  ��������l��$�0�������%0  u��������   ��������������  t[ǅ ���    �EP�˼����f��`�����`���Qh   ������R������P��������� ����� ��� t
ǅ����   �2�MQ������f��x����   k� ��x���������ǅ����   �������������J	  �EP�˖���������������� t�������y u#�p�������������P�������������e��������   t/�������B��������������+���������ǅ����   �(ǅ����    �������B��������������������  ������%0  u��������   �������������uǅX���������������X�����X����������MQ�˕������������������  ��   ������ u�t�������ǅ����   �������������������������������������������� t���������t��������������뾋�����+��������������u������ u�p��������������������������������������������������� t���������t��������������뾋�����+������������*  �MQ諔������D���膵������   3�tǅT���   �
ǅT���    ��T�����L�����L��� u&h�h�Yj h�  hx�j�o}������u̃�L��� uI�����    j h�  hx�h؛h�������ǅ���������� ����2����������	  �_  �������� t��D���f������f����D����������ǅ����   �%  ǅ����   �������� ��������������@������������������ǅ|���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Zh�  hp�j��������]  R�Bx���������������� t ��������������������]  ��|����
ǅ�����   �U���U�E�H��P��������������� ��������P������P������Q������R��|���P������Q������R�   k���0�R� �Ѓ�������%�   t6������ u-�� ����k���P������Q�   k�	��0�Q� �Ѓ���������gu:������%�   u-�� ����%���P������Q�   ����0�P� �Ѓ����������-u ������   ��������������������������R��������������  ��������@������ǅ����
   �   ǅ����
   �   ǅ����   ǅ����   �
ǅ����'   ǅ����   ��������   t2�   k� Ƅ����0��������Q�   �� ������ǅ����   �)ǅ����   ������%�   t��������   �������������� �  t�EP�������������������   ��������   t�UR�ƨ�����������������   �������� tE��������@t�UR�G���������������������EP�+���������������������@��������@t�UR���������������������EP������3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ������������������ }ǅ����   �%���������������������   ~
ǅ����   �����������u
ǅ����    �   i��  �������������������������������������������� �������������   �������RP������R������P�6�����0�������������RP������Q������R�r���������������������9~���������������������������������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0�������������������� �b  ��������@tv��������   t�   k� Ƅ����-ǅ����   �L��������t�   k� Ƅ����+ǅ����   �%��������t�   k� Ƅ���� ǅ����   ������+�����+�������l�����������u������Q�UR��l���Pj ��	  ����d���Q������R�EP������Q������R�"
  ����������t'��������u������R�EP��l���Qj0�	  �������� ��   ������ ��   ǅ<���    ��������t�����������h�����h�����������h�������h��������� ��   ��t���f�f��r�����r���Rj�E�P��4���Q聼������<�����t�������t�����<��� u	��4��� uǅ���������*��d���P������Q�UR��4���P�M�Q�	  ���N����(��d���R������P�MQ������R������P��  �������� |'��������t������R�EP��l���Qj �X  �������� tj������R�˂����ǅ����    ������������������ ��������������M�3�辒����]ÐW���ӡg�ʢ٢)���.�?���S�b� �I ��b�f�s��� ���ǤF����Ѩ�������e��+�ܮ   	
������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E����U�
�E��A��Q�]��������������������U��E����U�
�E��A�]�������U��E����U�
�E�f�A�]����������������������U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP葫�����E��}��u�M�������U����M���]�������������������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��|�U�    �E�E��M���M�}� ~N�U��E��MQ�UR�E�P�w������M���M�U�:�u�E�8*u�MQ�URj?�L�������띋E�8 u�M�U���]������������������������������������������������U��� �=� ��  �} t	�E�   ��E�    �E�E��}� u#hܥh�Yj jXh��j�mj������u̃}� u0记���    j jXh��h �hܥ�����������/  �} t	�E�   ��E�    �U�U�}� u#hx�h�Yj jYh��j��i������u̃}� u0�3����    j jYh��h �hx�萨���������   �M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���M�U���U�E���t�M��U�;��l����E��M�+���j �UR�EP��������]��������������������������������������������������������������������������������������������������������������������������������U���@�EP�M��3r���} t	�E�   ��E�    �M��M�}� u#hܥh�Yj j4h��j�.h������u̃}� u=�o����    j j4h��h�hܥ�̦�����E�����M�������E���  �} t	�E�   ��E�    �E�E�}� u#hx�h�Yj j5h��j�g������u̃}� u=�����    j j5h��h�hx��D������E�����M��u����E��;  �M��i�����   �����    ��   �M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���M�U���U�E���t�M��U�;��l����n�Ef�f�M��M�誳��P�U�R��c����f�E��E���E�Mf�f�U�M��}���P�E�P�c����f�E��M���M�U���t�E��M�;�t��U��E�+ЉUЍM��5����EЋ�]����������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P��SVW���1E�3�P�E�d�    �=� uEj�1f�����E�    �=� u�(  �������E������   �j�Z�����ËM�d�    Y_^[��]�������������������������������������������������U��j�h؊h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j�se�����E�    �EP�_   ���E��E������   �j訝����ËE�M�d�    Y_^[��]��������������������������������������������U����E�    j h9  h8�h��h���E�P�li����P�n�����}� u3��  �M�Q;|�u�E�H;����  �= � �G  �����uO���P���Q���R���Pj ���Q���R���P�M�QRjj�i  ��,�G���P���Q���R���P���Qj j ���R�E�HQj j�   ��,�l���uO�z�P�x�Q�v�R�t�Pj �p�Q�r�R�n�P�M�QRjj ��
  ��,�G�z�P�x�Q�v�R�t�P�r�Qj j �n�R�E�HQj j �
  ��,�   �E�   �E�   �E�   �E�   �U�zk}�E�   �E�   �E�
   �E�   j j j jj j �E�P�M�Q�U�BPjj�
  ��,j j j jj j �M�Q�U�R�E�HQjj ��	  ��,���;��}K�E�H;��|�U�B;��~3���   �M�Q;��~�E�H;��}
�   �   �F�U�B;��|�M�Q;��~
�   �   �E�H;��~�U�B;��}3��a�MkQ<�E�ʋUiB  �i��  �M�U�B;��u�M�;��|	�   ��3����U�;��}	�   ��3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���\~���M�]������������������U�������M�]������������������U���\����M�]������������������U��j�h��h�Ld�    P��SVW���1E�3�P�E�d�    j�J`�����E�    �J   �E������   �j艘����ËM�d�    Y_^[��]��������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    j�_�����E�    ������E�j h�   h8�h��h���E�P�f����P�,i����j h�   h8�h��h���M�Q��c����P�i����j h�   h8�h��h0��U�R蔁����P��h����轃���E�� �    �����������|�hh��������E�}� t�M������  �=� tj��P�Bl������    h(��@����=  � �   k(�<�M��n���tk|�<E��E������t$�=�� t�E�   ���+|�k�<�E���E�    �E�    �M�Qj j?�   k� �M܋Rj�h,�j �E�P� ��t"�}� u�   k� �   k�?�E܋� ��   k� �   k� �U܋
� �U�Rj j?�   �� �M܋Rj�h��j �E�P� ��t"�}� u�   �� �   k�?�U܋
� ��   �� �   k� �E܋� �E�   ��   �=� t"��P�M�Q蚆������u�E�   �   �=� tj��R�j����h  hl�j�E�P��������P��W�������=� u	�E�   �Aj h   h8�h��h���M�Q�U�R�ą������P��P������P�Kf�����M�Q�@������U�R�@������E�P�a������E������   �j蕔����Ã}� ��  j h3  h8�h��h��j�M�Qj@�   k� �M܋R������P��e�����E���E�M����-u�Eȃ��EȋM���M�U�R�;�����i�  �E��M����+t�E����0|�U����9�M���M��ԋU����:��   �M���M�U�R������k�<E��E��M����0|�E����9�U���U��ߋE����:u<�U���U�E�P蘟����E��E��M����0|�E����9�U���U��߃}� t�E��؉E��M����t	�E�   ��E�    �}� t@j hj  h8�h��hH�j�E�Pj@�   �� �U܋
P螥����P�^d������   �� �U܋
�  �M�Q�@������U�R�@������M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���VW�E�    �}�K  �E%  �yH���@��u�E��d   ����u#�El  ���  ����t�U�����E���M����U�E���E��M��Fi�m  M��E���������E����d   ��+��E+  ���  ����D1�   ���U��U�;U�E+E��M��k�U�ЉU���E+E�kMM�ȉM��}ud�U��  �yJ���B��u�E��d   ����u#�El  ���  ����t�U�����E���M����U��E�;E�~	�M����M��b�U��  �yJ���B��u�E��d   ����u#�El  ���  ����t�U�����E���M����U�E�E��M�M �M��}u2�U����kE$<E(k�<M,i��  U0����E�|��   �M����kU$<U(k�<E,i��  M0���j h�  h8�h��h0��U�R�!y����P�c`����iE��  �����y#����� \&������������*�=�� \&|���- \&������������U���_^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U�츜�]�������U�츠�]�������U�츘�]�������U��(�]�������U����} t	�E�   ��E�    �E��E��}� u#h�h�Yj j$hP�j��S������u̃}� u-�+����    j j$hP�h��h�舒�����   ��U����3���]���������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u#hؠh�Yj j-hP�j�*S������u̃}� u-�k����    j j-hP�h(�hؠ�ȑ�����   ��U����3���]���������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u#hH�h�Yj j6hP�j�jR������u̃}� u-諘���    j j6hP�hx�hH��������   ��U����3���]���������������������������������������������������U����} t�} w�} u�} t	�E�    ��E�   �E��E��}� u#h��h�Yj j?hP�j�Q������u̃}� u0�ٗ���    j j?hP�h`�h���6������   �_  �} t�   k� �M� �} t	�E�   ��E�    �U�U��}� u#h|�h�Yj jDhP�j�Q������u̃}� u0�I����    j jDhP�h`�h|�規�����   ��   �} t�}t	�E�    ��E�   �M�M�}� u#h��h�Yj jEhP�j�P������u̃}� u-�Ȗ���    j jEhP�h`�h���%������   �Q�E��(�Q�kz�������U��} u3��,�E�;Mv�"   ��U��(�P�MQ�UR舗������]�������������������������������������������������������������������������������������������������������������������������������������������U��Qh  �EP覄������u�M��_t	�E�    ��E�   �E���]�����������������������U��Qh  �EP�V�������u�M��_t	�E�    ��E�   �E���]�����������������������U����EP�M��X���M��ɛ����U���   �P�� �  �M��M��h���E���]�������������������������������U��h  �EP觃����]����������U��h  �EP臃����]����������U��Q�E��	u	�E�@   �j@�MQ�W������E��E���]������������������U��j �EP�*�����]�������������U��Qh  �EP��������u�M��_t	�E�    ��E�   �E���]�����������������������U��Qh  �EP趂������u�M��_t	�E�    ��E�   �E���]�����������������������U��j�EP�j�����]�������������U��h  �EP�G�����]����������U��j�EP�*�����]�������������U��hW  �EP������]����������U��j�EP������]�������������U��j�EP�ʁ����]�������������U��j�EP誁����]�������������U��h�   �EP臁����]����������U��j �EP�R�����]��������������U��h  �EP�G�����]����������U��h  �EP�'�����]����������U��Q�E=�   s	�E�   ��E�    �E���]�����������U��Q�E��	u	�E�@   �j@�MQ�ǀ�����E��E���]������������������U��j �EP蚀����]�������������U��j�EP�z�����]�������������U��h  �EP�W�����]����������U��j�EP�:�����]�������������U��hW  �EP������]����������U��j�EP������]�������������U��j�EP������]�������������U��j�EP�����]�������������U��h�   �EP�����]����������U��Q�E�    ��E����E��M���M�U�;Us�E���t�ڋE���]�����������������������U���  ���3ŉE��= � t3��M�3��h����]�� ��X  ����   Vh��� �5� ��tjh  ������QP�( ��tSh  ������P������P��  ����t4h 	  j ������P�օ���   �� ��Wujj ������P�օ�ugh 
  j h`��օ�uU�� ��WuHh  ������Pj �( ��t0h  ������P������P�C  ����tjj ������P�օ�u3�^�M�3��g����]�������������������������������������������������������������������������������������������U���$  ���3ŉE�S�� Wh   j hX��Ӌ���u,�� ��WuWWhX��Ӌ���u_3�[�M�3���f����]�V�5� hx�W�։�������tJh��W�։�������t8h��W�։�������t&������Pjj h��h  ���������tW�H^_3�[�M�3��\f����]Í�����ǅ����  P������P������Pj h ���������������������������W�H��u�������u���������u����r�If9�M�����x���f��M����\t�\   f��M����A���+����Q����A=  �C�������M��������M��������M��������M �������M���� ���M����$���M����(���M���f�,�h 	  f��M���������j P�Ӌ���u�� ��WujV������P�Ӌ��M���^_3�[�e����]������������������������������������������������������������������������������������������������������������������������������������������������������U���  ���3ŉE��E������V�uh   Qh   ������Qh   ������Qj�M�QP�fh����$��t3�^�M�3��d����]�hH�������j	P�S�������u�h<�������jP�9�������u�������P������P������P�E�P�uV�X���M������3�@^�c����]������������������������������������������������������������������U��E��D3��     �ES�]jf�K�E�PS�D��u3�[��]��u�u�u��( ��t�M��MZ  f9uًA<��~ҁ<PE  V�4t^3�[��]��F+��V��$�3�W3���t�;�r	��+�;X�rG��(;�r�;�t]G�=� u �=�� uJ����������t<������hx�P�� ��t�M�Qj j �M�Qj j j �u�Ѓ� ��u	_^3�[��]ËM�3ۉ]��=A�2�}  �M��U�Rh��S��P���c  �M�U�SSS�RVW�P ���B  �M�U��]�R��@h�Є��!  �M����  ��P����   �M��U�j R�U��R�UR�@�U�Rj �Є���   �E;�u�M�;�w	�E��;�r�M���P��u��   �E�����   =�����   ��Pj �(P�$�؅��}   �M��U�SRj ��U�j j R�@�Є�tP+u�;3rI�M��   ;�v
;4�r@;�r��D���U�M%��� j j j ��M�R�u��u܋@p�Є�t�E�   Sj �(P��M����]�M��P@�M��R8�M���R,_^��[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���<�} t�} v	�E�   ��E�    �E�E��}� u#hUh�Yj jh��j��@������u̃}� u0�%����    j jh��h�hU������   �  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R�Zg�����} t	�E�   ��E�    �E�E�}� u#h�Kh�Yj jh��j�@������u̃}� u0�G����    j jh��h�h�K�~�����   �  �U�U��E�E��}� v�M����t�E����E��M����M��܃}� ��   3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E��M���Qh�   �U��R�Lf��������t3�t	�E�   ��E�    �U܉U؃}� u#hP�h�Yj j h��j��>������u̃}� u0�2����    j j h��h�hP��}�����   �  �M��Uf�f��M���UċE����E��M���M�}� t�U����U�t�ƃ}� ��   3��Mf��}�tJ�}���tA�}v;�U��9h�s
�h��E��	�M���MԋU���Rh�   �E��P�.e����� L��t3�t	�E�   ��E�    �EЉẼ}� u#hPLh�Yj j*h��j��=������u̃}� u-����� "   j j*h��h�hPL�q|�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9h�s�h��U���E+E����M+ȉMȋU���Rh�   �E+E��M�TAR�?d����3���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���8�} u�} u�} u3��  �} t�} v	�E�   ��E�    �E�E��}� u#hUh�Yj jh��j�;������u̃}� u0������    j jh��h�hU�Yz�����   �  �} u`3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R�5b����3��&  �} ��   3��Mf��}�tJ�}���tA�}v;�U��9h�s
�h��E��	�M���M�U���Rh�   �E��P��a�����} t	�E�   ��E�    �M�M��}� u#h�Kh�Yj jh��j�x:������u̃}� u0蹀���    j jh��h�h�K�y�����   �I  �E�E��M�M��}�u?�U��Ef�f�
�U���E̋M����M��U���U�}� t�E����E�t���   �lo����t+�M;Mr#h Lh�Yj j+h��j�9������u̋E��Mf�f��E���MȋU����U��E���E�}� t�M����M�t�U���Ut뻃} u3��M�f��}� ��   �}�u3ҋE�Mf�TA��P   �J  3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E܋M���Qh�   �U��R��_����� L��t3�t	�E�   ��E�    �U؉Uԃ}� u#hPLh�Yj j>h��j�8������u̃}� u-��~��� "   j j>h��h�hPL�<w�����"   �r�}�tj�}���ta�M+M���;MsS�U+U����E+�9h�s�h��M���U+U����E+EЋM���Qh�   �U+U��E�LPQ�
_����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E�p�]����U����E�    �E�E��}� |,�}�~�}�t����M��U���~���E��t3�t	�E�   ��E�    �U�U��}� u#h,�h�Yj j?hp�j�M6������u̃}� u+�|���    j j?hp�hЦh,���t���������E���]�������������������������������������������������U���8�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E��}� u#hKh�Yj jh��j�{5������u̃}� u0�{���    j jh��h��hK�t�����   �v  �} u\�U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U�E�Ph�   �M��Q��[����3��  �} ��   �U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U�E�Ph�   �M��Q�[�����} t	�E�   ��E�    �U�U��}� u#h�Kh�Yj jh��j�?4������u̃}� u0�z���    j jh��h��h�K��r�����   �:  �M�M��U�U��}�u=�E��M���E���M̋U����U��E���E�}� t�M����M�t���   �5i����t+�U;Ur#h Lh�Yj j+h��j�3������u̋M��U���M���UȋE����E��M���M�}� t�U����U�t�E���Et뽃} u�M�� �}� ��   �}�u�UU�B� �P   �D  �E�  �}�tI�}���t@�}v:�M��9h�s�h��U��	�E���E܋M�Qh�   �U��R��Y����� L��t3�t	�E�   ��E�    �U؉Uԃ}� u#hPLh�Yj j>h��j�r2������u̃}� u-�x��� "   j j>h��h��hPL�q�����"   �p�}�th�}���t_�M+M���;MsQ�U+U����E+�9h�s�h��M���U+U����E+EЋM�Qh�   �U+U��E�LQ��X����3���]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    �E��Q�U�j j �EP�MQ�.�����E��}� u3���   �}� ~W3�uS�����3��u���rD�E���P�<������t#h��  �M��T	R�Z����P�r�����E���E�    �E��E���E�    �M�M��}� u3��u�U�R�E�P�MQ�UR�.������u�H�F�} uj j j j j��E�Pj �M�Q� �E��!j j �UR�EPj��M�Qj �U�R� �E�E�P�bG�����E��]����������������������������������������������������������������������������������������U����EP�M���8���MQ�UR�EP�MQ�M��)|��P�P������E��M��I���E���]����������������������������U����E�MH<�M��E�    �U��B�M��T�U���E���E�M���(�M��U��B9E�s#�M��U;Qr�E��H�U�J9Ms�E���3���]������������������������������U��j�h8�h�Ld�    P���SVW���1E�3�P�E�d�    �e��E�   �E�    �E�P�6^������u�E�    �E������E��   �M+M�MЋU�R�E�P�RZ�����E��}� u�E�    �E������E��}�M��Q$��   �u	�E�   ��E�    �E܉E��E������E��M�E������D�M���Eā}�  �u	�E�   ��E�    �E�Ëe��E�    �E������E���E������M�d�    Y_^[��]��������������������������������������������������������������������������������������U����E�E��M����MZ  t3��;�E��M�H<�M��U��:PE  t3�� �E����E�M����  t3���   ��]������������������������������������U��E��]����U���(V��P� �E��} t	�E�   ��E�    �M�M��}� u#h�h�Yj j>hH�j��+������u̃}� u0�+r���    j j>hH�h��h��j�����   ��  �E�     �}� ��  h   j hX��� �E��}� u�� ��Wuj j hX��� �E��}� uy3�t	�E�   ��E�    �U�U�}� u#h��h�Yj jVhH�j� +������u̃}� u0�aq���    j jVhH�h��h���i�����   ��   h,��M�Q�� �E��}� ��   3�t	�E�   ��E�    �E�E��}� u#h��h�Yj j\hH�j�*������u̃}� uD�� P�z\�������p���0j j\hH�h��h���i������ P�G\�����T�U�R� �E�j � �E؋Eܹ��;E�t
�U�R�Hj�EP�U���u�Jp���    �?p��� �3�^��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�} t,�}t&h�h�Yj h�   hH�j�)������u̋M�M��} tG�U��B%   t:�M�Q�Ul�����U��B%�����M��A�U��B    �E��     �M��A    ��]������������������������������������U����} u#ht�h�Yj j?hH�j�f(������u̋M�M��U�R��[����P�h������u3��  �`���    �� �9E�u	�E�    �#� `���    ���9E�u	�E�   �3���   �\����\��M��Q��  t3��   �E��<�� u\j[h��jh   ��#�����E�M��U����}� u0�E����E��M��U��Q�E��M���U��B   �E��@   �/�M��U�����A�M��U��B��M��A   �U��B   �E��H��  �U��J�   ��]�������������������������������������������������������������������������������������������������������U��3�]����������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E���M�����0��M��E�   �U�z uXj
�A'�����E�    �E�x u%j h�  �M��Q�T�����U�B���M�A�E������   �j
�W_����Ã}� t!�U���E������0��TR�  �E��M�d�    Y_^[��]��������������������������������������������������������������������U��j�hX�h�Ld�    P���SVW���1E�3�P�E�d�    �E������E�    j��o������u����:  j�&�����E�    �E�    �	�E����E��}�@��  �M��<�0� �  �U���0��E��	�M��@�M�U���0�   9E���   �M��Q����   �E�x uXj
�%�����E�   �M�y u%j h�  �U��R�S�����E�H���U�J�E�    �   �j
�]����Ã}� u+�E��P�  �M��Q��t�E��P� �=����}� u-�M��A�U�������E����M��U�+�0���E�������}��t��   ��   h�   h�jj@j �/<�����E�}� ��   �E��M��0��<��� �<��	�E��@�E�M���0���   9U�s#�E��@ �M�������U��B
�E��@    뿋M����M܋U����E܃�����0��D�U�R�Vn������u�E������������E������   �j�M\����ËE܋M�d�    Y_^[��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�} ��   �E;<���   �M���U������0��L����   �U���E������0��<�th�=p�u<�U�U��}� t�}�t�}�t�"j j��L�j j��L�
j j��L�E���M������0��
����3����g��� 	   �&���     �����]���������������������������������������������������������������U����}�u�K&���     �Eg��� 	   ����O  �} |�E;<�s	�E�   ��E�    �M��M��}� u&hMh�Yj h5  hP�j� ������u̃}� u<��%���     ��f��� 	   j h5  hP�h��hM�(_��������   �E���M������0��D
��t	�E�   ��E�    �M�M��}� u&h�Mh�Yj h6  hP�j��������u̃}� u9�0%���     �*f��� 	   j h6  hP�h��h�M�^���������E���M������0��
��]����������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E� �E��t
�M�� �M�U�� @  t�E��   �E�M��   t
�U���U�EP�� �E܃}� u�� P�h��������q  �}�u�M��@�M���}�u
�U���U��-:���E��}��u�d���    �#���     ����#  �E�    �EP�M�Q�=�����U���U�E����M�������0��E�D
�M����U�������0��L$�ဋU����E�������0��L$�E����M�������0��D
$$�M����U�������0��D$�E�   �E������   �K�}� u8�U����E�������0��T����E����M�������0��T�M�Q������Ã}� t�U��U���E������EԋM�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������U��Q�} ��   �E;<���   �M���U������0��<�um�=p�uB�M�M��}� t�}�t�}�t�(�URj��L��EPj��L��MQj��L�U���E������0��U�3����&b��� 	   �!���     �����]��������������������������������������������������������������U��E���M������0��D
P� ]�����������U����}�u�a��� 	   3��   �} |�E;<�s	�E�   ��E�    �M��M��}� u#hMh�Yj j(hةj��������u̃}� u*�(a��� 	   j j(hةh8�hM�Y����3���E���M������0��D
��@��]�������������������������������������������������U���,�} t�} u3��  �E���u�} t3ҋEf�3���  �MQ�M���#���M��'g����ztt3�M��g��� �xtt#hP�h�Yj jGhP�j��������u̍M���f����   �����    u*�} t�Mf��Ef��E�   �M��3���E��c  �M��f��P�M�R�g��������   �M��f��� �xt~\�M��of����U;Qt|J�} t	�E�   ��E�    �E�P�MQ�M��?f����BtP�MQj	�M��+f����BP� ��u?�M��f����U;Qtr�E�H��u"�7_��� *   �E������M���2���E��   �M���e����Bt�E�M���2���E��{�q�} t	�E�   ��E�    �M�Q�URj�EPj	�M��e����QR� ��u�^��� *   �E������M��a2���E���E�   �M��M2���E���M��@2����]����������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�[����]����������������������U��j�hȋh�Ld�    P���SVW���1E�3�P�E�d�    3�f�E�j�$�����E�    �MQ��\����f�E��E������   �j�WP�����f�E�M�d�    Y_^[��]������������������������������������������U��Q�=,��u����=,��u���  �(j �E�Pj�MQ�,�R�� ��u���  �f�E��]�����������������������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u�Z���     �T\��� 	   ����b  �} |�E;<�s	�E�   ��E�    �M��M܃}� u#hMh�Yj jTh��j�������u̃}� u9�����     ��[��� 	   j jTh��h�hM�=T���������  �E���M������0��D
��t	�E�   ��E�    �M؉Mԃ}� u#h�Mh�Yj jUh��j�������u̃}� u9�H���     �B[��� 	   j jUh��h�h�M�S��������5  �}���w	�E�   ��E�    �EЉẼ}� u#h$�h�Yj jVh��j�������u̃}� u9�����     �Z���    j jVh��h�h$��S��������   �UR�k_�����E�    �E���M������0��D
��t�MQ�UR�EP�4�����E��D�AZ��� 	   �1���     �E�����3�u#h(Nh�Yj jah��j�������u��E������   ��EP�a����ËE�M�d�    Y_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   V�E�    �E������E��p����}�u�����     ��X��� 	   �����  �} |�M;<�s	�E�   ��E�    �U��U��}� u&hMh�Yj h�   h��j�-������u̃}� u<�i���     �cX��� 	   j h�   h��hL�hM�P��������[  �M���U������0��L��t	�E�   ��E�    �U��U��}� u&h�Mh�Yj h�   h��j�������u̃}� u<�����     �W��� 	   j h�   h��hL�h�M�P��������  �}���w	�E�   ��E�    �M��M��}� u&h$�h�Yj h�   h��j��������u̃}� u<�8���     �2W���    j h�   h��hL�h$��O��������*  �E�    �} t �E���M������0��D
��t3���  �} tǅt���   �
ǅt���    ��t����M��}� u&hl�h�Yj h�   h��j�5������u̃}� u<�q���     �kV���    j h�   h��hL�hl���N��������c  �E���M������0��D
$�����E�M�M��}�t�}��&  �  �U��u	�E�   ��E�    �E��E��}� u&h`Qh�Yj h�   h��j�m������u̃}� u<����     �U���    j h�   h��hL�h`Q��M��������  �U���s	�E�   ��E��E��M��Mh�   h��j�UR������E�}� u�0U���    � ���    ����;  jj j �EP��5�����M���u������0��D1(�T1,�   �U��u	�E�   ��E�    �E��E��}� u&h`Qh�Yj h�   h��j�L������u̃}� u<����     �T���    j h�   h��hL�h`Q��L��������z  �U����U�E�E�M�MԋU���E������0��T��H��  �E���M������0��D
��
��  �} ��  �M���U������0��MԊT��Eԃ��EԋM���M�U���U�E���M������0��D

�E���?  �M���U������0�¹   k� �D%��
�  �} �  �M���U�����0��   k� �EԊL
%��Uԃ��UԋE���E�M���M�U���E�����0��   k� �D%
�E����   �M���U������0�¹   �� �T%��
tk�} te�E���M�����0��   �� �EԊL%��Uԃ��UԋE���E�M���M�U���E�����0��   �� �D%
�UR��K������tL�E���M������0��D
%�   t*��l���Q�U���E������0��R�� �E��}� tk�E��ubj �M�Q�U��R�E�P�M���U������0��Q�P��u!�� �E؋U�R�
�����E������
  �E����E��   j �M�Q�UR�E�P�M���U������0��Q�� ��t�}� |�U�;Uv^�� �E؃}�u#�.Q��� 	   ����M؉�E������
  �,�}�mu�E�    ��	  ��U�R�r	�����E�������	  �E�E܉E�M���U������0��L��   ��	  �U���  �}� tE�E����
u:�U���E������0��T���E���M������0��T�8�M���U������0��L����U���E������0��L�E�E��M��M��U�U�9U��?  �E������   �U���E������0��T��@u:�E���M������0��D
���M���U������0��D��U��E���
�U����U��E����E��  �  �M����t!�E��M����E����E��M����M��  �U�E�L�9M�sG�U��B��
u�M����M��U��
�E����E���M��U����M����M��U����U��)  �E����E��E�    j �M�Qj�U�R�E���M������0��
P�� ��u	�� �E؃}� u�}� u�M���U����U���   �E���M������0��D
��HtH�M��
u�U��
�E����E��,�M���U����U��E���M������0��E�D
�X�M�;M�u�U��
u�E�� 
�M����M��6jj�j��UR��.������x�����|����E��
t�M���U����U������E�+E�E��M���#  �}� �  �U����U��E����   u�U����U��e  �E�   �E����X���u"�}��E�;E�r�M����M��UЃ��U��͋E����X��U��}� u�0M��� *   �E������  �E���;E�u�M�MЉM���   �U���E������0��T��H��   �E���M������0��E�� �D
�M����M��}�|0�U���E�����0��   k� �M��	�L%�U����U��}�u0�E���M�����0��   �� �E�� �D%�M����M��U�+UЉU��"j�E��ؙRP�EP�-������x�����|����M�+M�M싕p�����R�EP�M�Q�U�Rj h��  � �E�}� u�� P�_�����E�������  �E�+E�9E�t	�E�   ��E�    �M���U������0��M��L0�U���U��  �}� �  �E�E��M��M�E�+����U�B9E���   �M����uB�E���M������0��D
���M���U������0��D�   �   �U����t �M��U�f�f��M����M��U���U��]�E�+����M�TA�9U�sI�E��H��
u�U���U��
   �M�f��U����U���E��M�f�f��E����E��M���M������U�+U�����U��l  �}� tE�E����
u:�U���E������0��T���E���M������0��T�8�M���U������0��L����U���E������0��L�E�E��M��M�U�U�9U���  �E������   �U���E������0��T��@u:�E���M������0��D
���M���U������0��D��U��E�f�f�
�U����U��E���E��9  �/  �M����t#�E��M�f�f��E����E��M���M��  �U�E�L�9M�sN�U��B��
u�M���M��
   �E�f��M����M���U��E�f�f�
�U����U��E���E��  �M���M��E�    j �U�Rj�E�P�M���U������0��Q�� ��u	�� �E؃}� u�}� u�   �E�f��M����M��6  �U���E������0��T��H��   �Ẽ�
u�
   �U�f�
�E����E��   �M̉Mĺ   �E�f��M����M��U���E������0��UĊ�T�Eă��EċM���U�����0��   k� �EĊ �D
%�M���U�����0��   �� �D%
�b�M�;M�u�Ũ�
u�
   �M�f��U����U��;jj�j��EP�)(������x�����|����M̃�
t�   �E�f��M����M��,����U�+U�U�E�;Et�M�Q��E�����}��u�U�U���EȉE��E�^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EP�MQ�UR�EP�����]��������������������U��EPj �MQh�l������]���������������������U���0�E�    3��EԉE؉E܉E��E�E�E�MЉM��} t	�E�   ��E�    �U��U�}� u&h��h�Yj h�  hЬj�#�������u̃}� u.�dA���    j h�  hЬhT�h���9��������C�M��A����U��BB   �E��@    �M��    �UR�EP�MQ�U�R�U���E��E���]��������������������������������������������������������������������U��EP�MQ�URh�l�_����]�������������������U��EPj �MQh�2�1����]���������������������U��EP�MQ�URh�2��
����]�������������������U��EPj �MQ�UR�����]����������������������U���H�E�    3��E��E��EĉEȉẺEЉEԍM��M��} t	�E�   ��E�    �U��U�}� u&h��h�Yj h�   hЬj�3�������u̃}� u1�t?���    j h�   hЬh4�h����7��������k  �} t	�E�   ��E�    �M��M�}� u&hX�h�Yj h�   hЬj��������u̃}� u1��>���    j h�   hЬh4�hX��O7���������   �E��@B   �M��U�Q�E��M��U��B����EP�MQ�UR�E�P�a?�����E��} u�E��   �M��Q���U�E��M�H�}� |"�U���  3Ɂ��   �M܋U�����M����U�Rj �+7�����E܋E��H���M�U��E�B�}� |!�M��� 3�%�   �E؋M�����E����M�Qj ��6�����E؋E���]�����������������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP�MQ������]��������������U���0�E������E�    �} t	�E�   ��E�    �E�E��}� u&h�h�Yj h9  hЬj�y�������u̃}� u1�<���    j h9  hЬh,�h��5��������9  �} u�} u�} u3��   �} t�} v	�E�   ��E�    �U�U�}� u&hحh�Yj h?  hЬj���������u̃}� u1�<���    j h?  hЬh,�hح�v4��������  �M;M��   ��;����U��EP�MQ�UR�E��P�MQh2�/*�����E��}����   �}�t^�}���tU�U��;UsJ�E���M+�9h�s�h��U���E���M+ȉM�U���Rh�   �E�M�TAR������@;���8"u
�6;���M�������  �c�";����U��EP�MQ�UR�EP�MQh2�u)�����E�3ҋE�Mf�TA��}��u"�}�u��:���8"u
��:���U������o  �}� ��   �   k� 3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E��M���Qh�   �U��R������}��u}3�t	�E�   ��E�    �M܉M؃}� u&h��h�Yj hf  hЬj���������u̃}� u1�:��� "   j hf  hЬh,�h���[2��������   ����{�}�t]�}���tT�E���;EsI�M����U+�9h�s
�h��E���M����U+щUԋE���Ph�   �M��U�DJP�0�����}� }	�E�������M��MЋEЋ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EPj �MQ�UR�EPh�l�&�����E��}� }	�E�������M��M��E���]�����������������������������U����EP�MQ�UR�EP�MQh�l�C&�����E��}� }	�E�������U��U��E���]���������������������������U���H�E�    3��E��E��EĉEȉẺEЉEԍM��M��} t	�E�   ��E�    �U�U��}� u&h��h�Yj h�   hЬj���������u̃}� u1�7���    j h�   hЬh��h���n/��������  �} t�} u	�E�    ��E�   �M�M�}� u&hP|h�Yj h�   hЬj�N�������u̃}� u1�6���    j h�   hЬh��hP|��.��������8  �E��@B   �M��U�Q�E��M��}���?v�U��B�����E���M��A�UR�EP�MQ�U�R�U���E��} u�E���   �}� ��   �E��H���M�U��E�B�}� |!�M��� 3�%�   �E��M�����E����M�Qj �.�����E��}��tY�U��B���E܋M��U܉Q�}� |"�E��� 3ҁ��   �U؋E�����U��
��E�Pj �T.�����E؃}��t�E�� 3ɋU�Ef�LP��M��y }�����������]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EPj �MQ�UR�EPh�2��"�����E��}� }	�E�������M��M��E���]�����������������������������U����EP�MQ�UR�EP�MQh�2�s"�����E��}� }	�E�������U��U��E���]���������������������������U���$�E������} t	�E�   ��E�    �E��E�}� u&h�h�Yj h  hЬj� �������u̃}� u1�a3���    j h  hЬh��h��+���������  �} t�} v	�E�   ��E�    �U��U�}� u&hحh�Yj h  hЬj��������u̃}� u1��2���    j h  hЬh��hح�6+��������x  �MQ�UR�EP�MQ�URh2�!�����E��}� }b�   k� 3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R�������}��uz3�t	�E�   ��E�    �M�M��}� u&h��h�Yj h  hЬj��������u̃}� u.��1��� "   j h  hЬh��h���'*��������l�}� |c�}�t]�}���tT�E���;EsI�M����U+�9h�s
�h��E���M����U+щU܋E���Ph�   �M��U�DJP�������E���]��������������������������������������������������������������������������������������������������������������������������������������������������������������������U��EPj �MQ�UR�EP������]������������������U����  ���3ŉE�ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    �EP��d����Y���ǅ����    ��/����P����} tǅH���   �
ǅH���    ��H�����L�����L��� u&h �h�Yj h  hx�j�-�������u̃�L��� uI�k/���    j h  hx�hT�h ���'����ǅ,���������d���������,����8  �} tǅ@���   �
ǅ@���    ��@�����8�����8��� u&h��h�Yj h  hx�j��������u̃�8��� uI��.���    j h  hx�hT�h���'����ǅ(���������d����G����(����  ǅ����    ǅ����    ǅ����    ǅ����    ǅt���    �Uf�f�������������� ����U���U�� ��� �  ������ �  �������� |%��������x�������������0����
ǅ0���    ��0���������������������������������������D�����D�����  ��D����$� Oǅ����   ������Q�UR������P�  ���J  ǅ����    ������������������������������������ǅ����    ǅ��������ǅ����    ��  �������������������� ������������wj��������8O�$� O���������������E���������������4���������������#�������ʀ   ����������������������e  ��������*u:�UR������������������� }���������������������ى������k�����
�������LЉ������  ǅ����    ��  ��������*u'�EP�t����������������� }
ǅ���������k�����
�������DЉ������  ��������������������I������������.�1  ��������`O�$�LO�U���lu�M���M��������   �����������������������   �M���6u+�E�H��4u�U���U������ �  �������   �M���3u(�E�H��2u�U���U������%����������S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    ������#�������� ���������������   �������D  ��������������������A������������7��
  ���������O�$��O��������0  u�������� ������ǅ����   �EP�m�����f�������������� ��   ���������   �   k� ������ǅT���   ��T���s��"����T���Ƅ���� ��d����B0��P��d����60��� �HtQ������R������P�5'������}
ǅ����   ��   k� f������f������������������ǅ����   �s	  �UR������������������ t�������x u#�p�������������R������������d������%   t/�������Q������������� �+���������ǅ����   �(ǅ����    �������Q���������������������  ��������0  u�������� �������������uǅ4���������������4�����4����������EP�������������������� ��   ������ u�p�������������������ǅ����    ���������������������;�����}O���������tB��d����X.��P�������P�e/������t������������������������������   ������ u�t�������ǅ����   ������������������������������������������ t���������t��������������뾋�����+��������������2  �UR�Q�������\����,������   3�tǅ`���   �
ǅ`���    ��`�����<�����<��� u&h�h�Yj h�  hx�j��������u̃�<��� uI�S&���    j h�  hx�hT�h������ǅ$���������d����������$���� 	  �g  �������� t��\���f������f����\����������ǅ����   �-  ǅ����   �������� f��������������@������������������ǅt���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Yh�  hp�j������]  P������������������� t ��������������������]  ��t����
ǅ�����   �E���E�M�Q��A�������������d����x+��P������Q������R������P��t���Q������R�����P�   k���0�P� �Ѓ���������   t6������ u-��d����+��P������R�   k�	��0�R� �Ѓ���������gu;��������   u-��d�����*��P������R�   ����0�Q� �Ѓ����������-u!��������   ��������������������������P�������������  ��������@������ǅ����
   �   ǅ����
   �   ǅ����   ǅ����   �
ǅ����'   ǅ����   ��������   t8�   k� �0   f��������������Q�   �� f������ǅ����   �)ǅ����   ��������   t������   �������������� �  t�UR������������������   ������%   t�MQ�d�����������������   �������� tE��������@t�MQ�����������������������UR�����������������������@��������@t�MQ���������������������UR������3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ������������������ }ǅ����   �%���������������������   ~
ǅ����   �����������u
ǅ����    �   i��  ������������������������������������������ �������������   �������RP������R������P�������0�������������RP������Q������R����������������������9~���������������������������������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0�������������������� �a  ��������@��   ��������   t!�   k� �-   f������ǅ����   �V��������t!�   k� �+   f������ǅ����   �*��������t�   k� �    f������ǅ����   ������+�����+�������|�����������u������Q�UR��|���Pj �  ����P���Q������R�EP������Q������R�  ����������t'��������u������R�EP��|���Qj0�;  �������� ��   ������ ��   ��������������������x�����x����������x�������x�������� ��   ��d�����$��P��d����$��� �HtQ������R������P�������X�����X��� ǅ���������2������Q�UR������P��  ���������X����������X����(��P���R������P�MQ������R������P�  �������� |'��������t������R�EP��|���Qj �  �������� tj������R�j�����ǅ����    ������������������d�������������M�3��]�����]�\>�>�>k?�?�?-@�A2?C?!??W?f? �I �@dAj@uA�A �F�A~C|H�B,F�AEHE�HrH�CcH�H>L   	
����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E�H��@t�U�z u�E����U�
�4�EP�MQ������Ё���  u�E� ������M����E�]�������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�U������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��~�U�    �E�E��M���M�}� ~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������뛋E�8 u�M�U���]����������������������������������������������U���<�} t�} v	�E�   ��E�    �E�E��}� u#hKh�Yj jh��j�d�������u̃}� u0����    j jh��hp�hK������   �o  �} ��   �U� �}�tI�}���t@�}v:�E��9h�s�h��M��	�U���U�E�Ph�   �M��Q��������} t	�E�   ��E�    �U�U�}� u#h�Kh�Yj jh��j��������u̃}� u0�����    j jh��hp�h�K�(�����   �  �M�M��U�U��}� v�E����t�U����U��E����E��܃}� ��   �M� �}�tH�}���t?�}v9�U��9h�s
�h��E��	�M���M��U�Rh�   �E��P�����������t3�t	�E�   ��E�    �E܉E؃}� u#hP�h�Yj j h��j�z�������u̃}� u0����    j j h��hp�hP�������   �  �U��E��
�U���EċM����M��U���U�}� t�E����E�t�ȃ}� ��   �M� �}�tH�}���t?�}v9�U��9h�s
�h��E��	�M���MԋU�Rh�   �E��P������� L��t3�t	�E�   ��E�    �EЉẼ}� u#hPLh�Yj j*h��j�b�������u̃}� u-���� "   j j*h��hp�hPL� 
�����"   �p�}�th�}���t_�U+U���;UsQ�E+E����M+�9h�s�h��U���E+E����M+ȉMȋU�Rh�   �E+E��M�TR�������3���]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���L�U�M�}� t	�E�   ��E�    �E��E܃}� u&h�uh�Yj h>  h��j�a�������u̃}� u3����    j h>  h��h��h�u�������   �  �}� v	�E�   ��E�    �U؉Uԃ}� u&h��h�Yj h?  h��j���������u̃}� u3�!���    j h?  h��h��h���{�����   �  �M�� �}��tH�}����t?�}�v9�U��9h�s
�h��E��	�M���MЋU�Rh�   �E��P�b������} t	�E�   ��E�   �M�;M�v	�E�   ��E�    �UȉUă}� u&h �h�Yj hA  h��j���������u̃}� u3�4��� "   j hA  h��h��h �������"   �)  �}r�}$w	�E�   ��E�    �M��M��}� u&h��h�Yj hB  h��j�l�������u̃}� u3����    j hB  h��h��h��������   �  �E�    �E�E��} t+�M��-�U����U��E����E��M�ًU�� �ډM�U�E��E�M3�RQ�EP�MQ�h����E�U3�PR�MQ�UR�����E�U�}�	v�E��W�M���U����U���E��0�M���U����U��E����E��} w�} v�M�;M�r��U�;U���   �   k� �U��
 �E�;E�s	�E�   ��E�    �M��M��}� u&h��h�Yj hf  h��j��������u̃}� u0�M��� "   j hf  h��h��h��������"   �E�E��  �M����M��U���E��M��U���M�U���E����E��M���M�U�;U�r�3���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�}�����]��������������������������U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP��   �E��j �MQ�UR�EP�MQ��   �E��E���]�����������������������������U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ�w   ��]��������������������U��j �EP�MQ�UR�U�M����]�������������������U��j �EP�MQ�UR�EP�   ]���������������������U���D�} t	�E�   ��E�    �E�E�}� u#h�uh�Yj jfh��j��������u̃}� u0�����    j jfh��h�h�u�H�����   �Y  �} v	�E�   ��E�    �U��U܃}� u#h��h�Yj jgh��j�/�������u̃}� u0�p���    j jgh��h�h���� �����   ��  �M� �}�tH�}���t?�}v9�U��9h�s
�h��E��	�M���M؋U�Rh�   �E��P�������} t	�E�   ��E�   �M;M�v	�E�   ��E�    �UЉŨ}� u#h �h�Yj jih��j�H�������u̃}� u0���� "   j jih��h�h ���������"   ��  �}r�}$w	�E�   ��E�    �MȉMă}� u#h��h�Yj jjh��j���������u̃}� u0����    j jjh��h�h���e������   �v  �E�    �E�E��} t �M��-�U����U��E���E�M�ىM�U��U��E3��u�U�E3��u�E�}�	v�E��W�M���U����U���E��0�M���U����U��E���E�} v�M�;Mr��U�;U��   �   k� �U�
 �E�;Es	�E�   ��E�    �M��M��}� u&h��h�Yj h�   h��j薿������u̃}� u0����� "   j h�   h��h�h���1������"   �E�E��  �M����M��U���E��M��U����M��U���E����E��M����M��U�;U�r�3���]� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���L�U�M�}� t	�E�   ��E�    �E��E܃}� u&h�uh�Yj h>  h��j���������u̃}� u3����    j h>  h��h�h�u�\������   �  �}� v	�E�   ��E�    �U؉Uԃ}� u&h��h�Yj h?  h��j�@�������u̃}� u3����    j h?  h��h�h����������   �,  3ɋU�f�
�}��tK�}����tB�}�v<�E��9h�s�h��M��	�U���UЋE���Ph�   �M��Q�������} t	�E�   ��E�   �U�;U�v	�E�   ��E�    �EȉEă}� u&h �h�Yj hA  h��j�N�������u̃}� u3���� "   j hA  h��h�h ���������"   �:  �}r�}$w	�E�   ��E�    �U��U��}� u&h��h�Yj hB  h��j�ǻ������u̃}� u3����    j hB  h��h�h���b������   �  �E�    �M�M��} t0�-   �E�f��M����M��U����U��E�؋M�� �ىE�M�U��U�E3�QP�UR�EP�����E�M3�RQ�EP�MQ�����E�U�}�	v�U��W�E�f��M����M���U��0�E�f��M����M��U����U��} w�} v�E�;E�r��M�;M���   �   k� 3ɋU�f��E�;E�s	�E�   ��E�    �M��M��}� u&h��h�Yj hf  h��j�^�������u̃}� u0� ��� "   j hf  h��h�h����������"   �M3��M�f��U����U��E�f�f�M��U��E�f�f�
�U�f�E�f��M����M��U���U�E�;E�r�3���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�}
u�} |�} s	�E�   ��E�    �E�P�MQ�UR�EP�U�M�m�����]��������������������������U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP��   �E��j �MQ�UR�EP�MQ��   �E��E���]�����������������������������U��Q�}
u�} }	�E�   ��E�    �E�P�MQ�UR�EP�MQ�w   ��]��������������������U��j �EP�MQ�UR�U�M�t���]�������������������U��j �EP�MQ�UR�EP�   ]���������������������U���D�} t	�E�   ��E�    �E�E�}� u#h�uh�Yj jfh��j���������u̃}� u0�;����    j jfh��h�h�u�������   �o  �} v	�E�   ��E�    �U��U܃}� u#h��h�Yj jgh��j��������u̃}� u0������    j jgh��h�h���������   ��  3ɋUf�
�}�tK�}���tB�}v<�E��9h�s�h��M��	�U���U؋E���Ph�   �M��Q��������} t	�E�   ��E�   �U;U�v	�E�   ��E�    �EЉẼ}� u#h �h�Yj jih��j蓵������u̃}� u0������ "   j jih��h�h ��1������"   �  �}r�}$w	�E�   ��E�    �UȉUă}� u#h��h�Yj jjh��j��������u̃}� u0�S����    j jjh��h�h���������   �  �E�    �M�M��} t%�-   �E�f��M����M��U���U�E�؉E�M��M��E3��u�U�E3��u�E�}�	v�U��W�E�f��M����M���U��0�E�f��M����M��U���U�} v�E�;Er��M�;M��   �   k� 3ɋUf��E�;Es	�E�   ��E�    �M��M��}� u&h��h�Yj h�   h��j�س������u̃}� u0����� "   j h�   h��h�h���s������"   �M3��M�f��U����U��E�f�f�M��U��E�f�f�
�U�f�E�f��M����M��U����U��E�;E�r�3���]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��} u�  �E�H;4�tj�U�BP�������M�Q;8�tj�E�HQ�������U�B;<�tj�M�QR�u������E�H;@�tj�U�BP�V������M�Q;D�tj�E�HQ�7������U�B ;H�tj�M�Q R�������E�H$;L�tj�U�B$P��������M�Q8;`�tj�E�H8Q�ڿ�����U�B<;d�tj�M�Q<R軿�����E�H@;h�tj�U�B@P蜿�����M�QD;l�tj�E�HDQ�}������U�BH;p�tj�M�QHR�^������E�HL;t�tj�U�BLP�?�����]��������������������������������������������������������������������������������������������������������������U���VW�E�    �E�E��E�    �   k��E���    u�   ���U��
�    �n  jSh4�jjPj�D������E��}� u
�   �  jYh4�jj�̫�����E�}� uj�E�P�4������   ��  �M��    �   k��M���    �o  jeh4�jj�v������E��}� u&j�U�R�޽����j�E�P�н�����   �u  �M��    �   k��M���   �U��E�    �E���Pj�M�Qj�U�R�K�����E��E��E���Pj�M�Qj�U�R�*�����E��E��E���Pj�M�Qj�U�R�	�����E��E��E���Pj�M�Qj�U�R�������E��E��E���Pj�M�Qj�U�R�������E��E��E��� PjP�M�Qj�U�R������E��E��E���$PjQ�M�Qj�U�R������E��E��E���(Pj�M�Qj �U�R�d�����E��E��E���)Pj�M�Qj �U�R�C�����E��E��E���*PjT�M�Qj �U�R�"�����E��E��E���+PjU�M�Qj �U�R������E��E��E���,PjV�M�Qj �U�R�������E��E��E���-PjW�M�Qj �U�R������E��E��E���.PjR�M�Qj �U�R������E��E��E���/PjS�M�Qj �U�R�}�����E��E��E���8Pj�M�Qj�U�R�\�����E��E��E���<Pj�M�Qj�U�R�;�����E��E��E���@Pj�M�Qj�U�R������E��E��E���DPj�M�Qj�U�R�������E��E��E���HPjP�M�Qj�U�R�������E��E��E���LPjQ�M�Qj�U�R������E��E�t@�E�P������j�M�Q�к����j�U�R�º����j�E�P贺�����   �Y  �M��QR�  ����   �(��}��E���   �U����M���   �E��J�H�U���   �M��P�Q�E���   �U��A0�B0�M���   �E��J4�H4�U��   �}� t	�E��    ��E�    �E�    �E�(��M���    tE�U���   �����Iu2�U���    w&hd�h�Yj h�   h��j��������u̋M�yx t5�U�Bx�����Iu%j�U���   P腹����j�M�QxR�t������E�M����   �U�E�Bx�M�U����   3�_^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]������������������������������������U��} u�   �E�;(�tj�U�P�������M�Q;,�tj�E�HQ��������U�B;0�tj�M�QR�׶�����E�H0;X�tj�U�B0P踶�����M�Q4;\�tj�E�H4Q虶����]��������������������������������������������������������U���VW�E�    �E�    �E�E��E�    �   ���U��
�    u�   k��U��
�    �1  jeh�jjPj�Ϳ�����E��}� u
�   ��  �E�   ���   �}��jqh�jj�B������E��}� uj�M�Q誵�����   �}  �U��    �   ���M���    �E  j}h�jj�������E�}� u&j�U�R�T�����j�E�P�F������   �  �M��    �   ���E���   �M�U�Rj�E�Pj�M�Q�������E��E��U���Rj�E�Pj�M�Q������E��E��U���Rj�E�Pj�M�Q������E��E��U���0Rj�E�Pj�M�Q�h�����E��E��U���4Rj�E�Pj�M�Q�G�����E��E�t0�U�R�K�����j�E�P�`�����j�M�Q�R���������'  �U��BP��  ���A�E�    �M��(���E��,��H�U��0��B�M��X��Q0�E��\��H4�U��   �}� t	�E��    ��E�    �E�    �E�(��M�y| t?�U�B|�����Iu/�U�z| w&h@�h�Yj h�   h��j��������u̋M�yx t5�U�Bx�����Iu%j�U�BxP�W�����j�M���   R�C������E�M�H|�U�E��Bx�M�U����   3�_^��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E���tk�U���0|$�M���9�E���0�U�
�E���E�:�M���;u&�E�E��M��U��B��M����M��U����u��	�M���M닋�]������������������������������������U��} u�	  j�   �� �M�R�y�����j�   ���M�R�a�����j�   k��U�
P�H�����j�   ���U�
P�/�����j�   k��E�Q������j�   k��M�R�������j�   k� �U�
P������j�   �� �U�D
P�ʰ����j�   ��U�D
P豰����j�   k��E�LQ藰����j�   ���E�LQ�}�����j�   k��M�TR�c�����j�   k��U�D
P�I�����j�   k� �E�LQ�/�����j�   k� �M�T8R������j�   �� �M�T8R�������j�   ���M�T8R������j�   k��U�D
8P�ȯ����j�   ���U�D
8P讯����j�   k��E�L8Q蔯����j�   k��M�T8R�z�����j�   k��U�D
8P�`�����j�   ���U�D
8P�F�����j�   k�	�E�L8Q�,�����j�   k�
�M�T8R������j�   k��U�D
8P�������j�   k� �E�LhQ�ޮ����j�   �� �E�LhQ�Į����j�   ��E�LhQ諮����j�   k��M�ThR葮����j�   ���M�ThR�w�����j�   k��U�D
hP�]�����j�   k��E�LhQ�C�����j�   k��M�ThR�)�����j�   ���M�ThR������j�   k�	�U�D
hP�������j�   k�
�E�LhQ�ۭ����j�   k��M�ThR�������j�   k� �U��
�   P褭����j�   �� �U��
�   P臭����j�M���   R�s�����j�E���   Q�_�����j�U���   P�K�����j�   �� �U��
�   P�.�����j�   ��U��
�   P������j�   k��E���   Q�������j�   ���E���   Q�ج����j�   k��M���   R軬����j�   k��U��
�   P螬����j�   k� �E���   Q聬����j�   �� �E���   Q�d�����j�   ��E���   Q�H�����j�   k��M���   R�+�����j�   ���M���   R������j�   k��U��
�   P������j�   k��E���   Q�ԫ����j�   k� �M���   R跫����j�   k� �U��
�   P蚫����j�   �� �U��
�   P�}�����j�   ��U��
�   P�a�����j�   k��E���   Q�D�����j�   ���E���   Q�'�����j�   k��M���   R�
�����j�   k��U��
�   P������j�   k��E���   Q�Ъ����j�   ���E���   Q質����j�   k�	�M���   R薪����j�   k�
�U��
�   P�y�����j�   k��E���   Q�\�����j�   k� �M��  R�?�����j�   �� �M��  R�"�����j�   ���M��  R������j�   k��U��
  P������j�   ���U��
  P�̩����j�   k��E��  Q诩����j�   k��M��  R蒩����j�   k��U��
  P�u�����j�   ���U��
  P�X�����j�   k�	�E��  Q�;�����j�   k�
�M��  R������j�   k��U��
  P������j�   k� �E��L  Q������j�   �� �E��L  Q�Ǩ����j�U��T  P賨����j�M��X  R蟨����j�E��\  Q苨����j�U��`  P�w�����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�   k��U��
�    trj@h�jhd  j�¯�����E��}� u
�   �   �EP�M�Q��   ����t$�U�R�������j�E�P讥�����   �   �M�ǁ�      ��E����U���   ��tN�E���   ���   �����Ju5�E���   ���    #h �h�Yj jPhx�j薖������u̋E�M����   3���]��������������������������������������������������������������������������������U����E�    �   k��U��
�   �E��   k��E���   �M�} u����  �U�R艽�����M��`  �U�U��E�    �   �� EPj1�M�Qj�U�R������E��E��   ��EPj2�M�Qj�U�R�������E��E��   k�MQj3�U�Rj�E�P�������E��E��   ��MQj4�U�Rj�E�P������E��E��   k�URj5�E�Pj�M�Q�w�����E��E��   k�EPj6�M�Qj�U�R�Q�����E��E��   k� MQj7�U�Rj�E�P�+�����E��E��   �� �U�D
Pj*�M�Qj�U�R������E��E��   ���M�TRj+�E�Pj�M�Q�ؿ����E��E��   k��M�TRj,�E�Pj�M�Q访����E��E��   ���E�LQj-�U�Rj�E�P脿����E��E��   k��E�LQj.�U�Rj�E�P�Z�����E��E��   k��E�LQj/�U�Rj�E�P�0�����E��E��   k� �E�LQj0�U�Rj�E�P������E��E��   k� �E�L8QjD�U�Rj�E�P�ܾ����E��E��   �� �U�D
8PjE�M�Qj�U�R貾����E��E��   ���M�T8RjF�E�Pj�M�Q艾����E��E��   k��M�T8RjG�E�Pj�M�Q�_�����E��E��   ���E�L8QjH�U�Rj�E�P�5�����E��E��   k��E�L8QjI�U�Rj�E�P������E��E��   k��E�L8QjJ�U�Rj�E�P������E��E��   k��E�L8QjK�U�Rj�E�P跽����E��E��   ���U�D
8PjL�M�Qj�U�R荽����E��E��   k�	�U�D
8PjM�M�Qj�U�R�c�����E��E��   k�
�U�D
8PjN�M�Qj�U�R�9�����E��E��   k��U�D
8PjO�M�Qj�U�R������E��E��   k� �U�D
hPj8�M�Qj�U�R������E��E��   �� �M�ThRj9�E�Pj�M�Q軼����E��E��   ��E�LhQj:�U�Rj�E�P蒼����E��E��   k��E�LhQj;�U�Rj�E�P�h�����E��E��   ���U�D
hPj<�M�Qj�U�R�>�����E��E��   k��U�D
hPj=�M�Qj�U�R������E��E��   k��U�D
hPj>�M�Qj�U�R������E��E��   k��U�D
hPj?�M�Qj�U�R�������E��E��   ���M�ThRj@�E�Pj�M�Q薻����E��E��   k�	�M�ThRjA�E�Pj�M�Q�l�����E��E��   k�
�M�ThRjB�E�Pj�M�Q�B�����E��E��   k��M�ThRjC�E�Pj�M�Q������E��E��   k� �M���   Rj(�E�Pj�M�Q������E��E��   �� �E���   Qj)�U�Rj�E�P辺����E��E��M���   Qj�U�Rj�E�P蚺����E��E��M���   Qj �U�Rj�E�P�v�����E��E��M���   Qh  �U�Rj�E�P�O�����E��E��M���   Qh	  �U�Rj �E�P�(�����E��E��   �� �U��
�   Pj1�M�Qj�U�R�������E��E��   ���M���   Rj2�E�Pj�M�Q�Ϲ����E��E��   k��M���   Rj3�E�Pj�M�Q袹����E��E��   ���E���   Qj4�U�Rj�E�P�u�����E��E��   k��E���   Qj5�U�Rj�E�P�H�����E��E��   k��E���   Qj6�U�Rj�E�P������E��E��   k� �E���   Qj7�U�Rj�E�P������E��E��   �� �U��
�   Pj*�M�Qj�U�R�������E��E��   ���M���   Rj+�E�Pj�M�Q蕸����E��E��   k��M���   Rj,�E�Pj�M�Q�h�����E��E��   ���E���   Qj-�U�Rj�E�P�;�����E��E��   k��E���   Qj.�U�Rj�E�P������E��E��   k��E���   Qj/�U�Rj�E�P������E��E��   k� �E���   Qj0�U�Rj�E�P贷����E��E��   k� �E���   QjD�U�Rj�E�P臷����E��E��   �� �U��
�   PjE�M�Qj�U�R�Z�����E��E��   ���M���   RjF�E�Pj�M�Q�.�����E��E��   k��M���   RjG�E�Pj�M�Q������E��E��   ���E���   QjH�U�Rj�E�P�Զ����E��E��   k��E���   QjI�U�Rj�E�P觶����E��E��   k��E���   QjJ�U�Rj�E�P�z�����E��E��   k��E���   QjK�U�Rj�E�P�M�����E��E��   ���U��
�   PjL�M�Qj�U�R� �����E��E��   k�	�U��
�   PjM�M�Qj�U�R������E��E��   k�
�U��
�   PjN�M�Qj�U�R�Ƶ����E��E��   k��U��
�   PjO�M�Qj�U�R虵����E��E��   k� �U��
  Pj8�M�Qj�U�R�l�����E��E��   �� �M��  Rj9�E�Pj�M�Q�?�����E��E��   ��E��  Qj:�U�Rj�E�P������E��E��   k��E��  Qj;�U�Rj�E�P������E��E��   ���U��
  Pj<�M�Qj�U�R蹴����E��E��   k��U��
  Pj=�M�Qj�U�R茴����E��E��   k��U��
  Pj>�M�Qj�U�R�_�����E��E��   k��U��
  Pj?�M�Qj�U�R�2�����E��E��   ���M��  Rj@�E�Pj�M�Q������E��E��   k�	�M��  RjA�E�Pj�M�Q�س����E��E��   k�
�M��  RjB�E�Pj�M�Q諳����E��E��   k��M��  RjC�E�Pj�M�Q�~�����E��E��   k� �M��L  Rj(�E�Pj�M�Q�Q�����E��E��   �� �E��L  Qj)�U�Rj�E�P�$�����E��E��M��T  Qj�U�Rj�E�P� �����E��E��M��X  Qj �U�Rj�E�P�ܲ����E��E��M��\  Qh  �U�Rj�E�P赲����E��E��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��SVWUj j h(��u胹��]_^[��]ËL$�A   �   t2�D$�H�3��	���U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h0�d�5    ���3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y0�u�Q�R9Qu�   �SQ����SQ����L$�K�C�kUQPXY]Y[� ��������������������������������������������������������������������������������������������U��Q�M��E��     �E���]����������U����M��E��H�� ����U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M�9 ��  �U������  �E�    �U��E���M����E��M�����  �M���M;���   �U����_��   �U����$��   �U����<��   �U����>��   �U����-tw�U����a|�U����z~]�U����A|�U����Z~C�U����0|�U����9~)�U�����   |�U�����   ~	�tz����t�U����U���E��H�� ������U��J�   ������E�P�M�Q�M��v����U����tG�U���M��U�U�E����U�
�E�;E�t�M��Q�� ������E��P�M��    � �M��6�����u�U��B% ������M��A��U��B% ������M��A��U��B% ������M��A�E���]� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M��E��M���I�H�E���]� ����������������U��Q�M��E��H�� ����U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M��"����E���]� ���������������������������������������������������������������U����M��} tpj h@�j�މ�����E��}� t�EP�M��e����E���E�    �M��U��E��8 t	�E�    ��E�   �M����   �U��B% �����M��A��U��B% ����M��A�U��    �E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E���]� ������������������������������������������������������������������������������U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} t%�MQ�m�  ���E��}� v�U�R�EP�M��{����E���]� ������������������������������������������������������������������������U����M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�}t�}t	�E�    ��E�E��M����   �U��B% �����M��A�U��    �}u.�EP�m������M���U��: u�E��H�� ������U��J�E���]� ��������������������������������������������������������������������������U��Q�M��E��     �M��Q�� ����E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�E���]��������������������������������������������������������U���(���3ŉE��M��E��E؋M��Q�� ����E��P�M��    �U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%����M��A�U�� �E� �} |�} s�E��E�؋M�� �ىE�M�U؃��U�j j
�EP�MQ譐����0�� �U؈j j
�EP�MQ�����E�U�UUu��E߅�t�M؃��M؋U��-�E؍M�+��   +�R�E�P�M��x����E��M�3��z�����]� �����������������������������������������������������������������������������������������������������������U���$���3ŉE��M��E��E܋M��Q�� ����E��P�M��    �U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%�����M��A�U��B%����M��A�U�� �E܃��E�j j
�MQ�UR�������0�� �M܈j j
�UR�EP�;����E�U�MMu��U܍E�+й   +�Q�U�R�M��ج���E��M�3��ړ����]� �������������������������������������������������������������������������������������������U��Q�M��E�� ��E���]����������U����M��M�輈���E�� l��M��U�Q�E��xu	�E�   ��E�    �M��U��Q�E���]� ����������������������������������U��Q�M��E�� �����E���]����������U��Q�M��M�������M���,赹���E�(��(��$��} t�U�0��E�,���,�    �0�    �M���,���U����E�4��M�<��8� �E���]� �����������������������������������������������U��Q�M��M��n����E�� 0��M��U�Q�E���]� ����������������������U����M��M��,����E�� X��} t#�M譙����t�M蠙����u	�E�    ��M�M��U��E��B�E���]� �������������������������������������U��Q�M��M�讆���E�� ���M��U�Q�E��M�H�U��B�����E���]� �������������������U����M��M��\����E�� D��} t\�} tVj h@��MQ��~�����E��U��E��B�M��U�Q�E��x t�MQ�UR�E��HQ��  ���
�U��B    ��E��@    �M��A    �E���]� ���������������������������������������U��EP�MQ�@�����]����������U��Q�M��E��M���I�H�E���]� ����������������U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�M��tj�UR�M������E���]� ���������������������������������������������������������������U����M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�} tXj h@�j�#|�����E��}� t�MQ�M�誖���E���E�    �U��E��M��9 u�U��B% ������M��A��U��B% ������M��A�E���]� ���������������������������������������������������������������������������������U��Q�M��E��H�� ����U��J�E��     �M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q�������E��P�M��Q������E��P�MQ�e�  ��P�UR�M������E���]� ������������������������������������������������������������U��Q�M��E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H�������U��J�E��H������U��J�E%�   �M��Q�� ���ЋE��P�}u0�MQ裃�����U���E��8 u�M��Q�� ������E��P�	�M��    �E���]� ���������������������������������������������������������������������U��Q�M��} |�}	~j�M�:����E�;�9�E��8�t
�M��U;~j�M�����E���E�M��T�R�M��w���E��]� �����������������������������U���H�M��M�������M�������=(� �E  �(����?uQ�   �� �(����@u;�$����$��E�P�op����PhL��M�Q��z����P�M��f����   �(����?ut�   �� �(��
��$u]j �M�Q��}����P�M��tf���M��͑����t��}����u.�$����t!�(��$��U�R��o����P�M��0f���e�   k� �(��
��?u9�   �� �(��
��?u"�   ��(��
��@uj�M�萍����M�Q�qo����P�M���e���M��"�����u	3��  �@�M�������t�4}����u�$����t�(�Q�M��ɚ����U�R�M��se���=,� u1�M�辮�����0�jh@��0�P�v�����E�M�,��=,� ��   �0�R�,�P�M��ڦ���,��M��U��U��E����tY�U���� u0�M����M��U�� �E����E��M���� u�E����E�����M��U����M����M��U����U�띋E��M����,���]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EP�MQ�UR�M��2����������E��]������������������������U����EP�MQ�UR�M�肱�����Ҍ���E��]�������������������������U����EP�MQ�UR�M�������蒌���E��]�������������������������U����M��E�P�M��s���MQ�M�������U�R�M�ss���E��]� ��������������������������U����M��E�P�M��;s���MQ�M��h����U�R�M�"s���E��]� �������������������������U����M��E�P�M���r���MQ�M��ӫ���U�R�M��r���E��]� ��������������������������U����M��E�P�M��r���MQ�M��u����U�R�M�r���E��]� ��������������������������U����M��E�P�M��Kr���MQ�M��ͱ���U�R�M�3r���E��]� ��������������������������U��Q�M��M��n����tG�M�o����t�M�Ό��P�M��n����(�M���n����t�EP�M��Ja����M�R�M��>v���E���]� �����������������������������U����M��M��n����tb�E��tZ�M��n����t�MQ�M��Dx���?j h@�j�5r�����E��}� t�UR�M�������E���E�    �E�P�M��u���E���]� ��������������������������������U����M��M��tm������   �} ��   �M���m����t�EP�M���f���j�M萋����t�M脋����u@j h@�j�wq�����E��}� t�MQ�M�������E���E�    �U�R�M���t����M�7���P�M��ׯ���E���]� ������������������������������������������������U����M��M��l����tu�} to�E���te�M��	m����t�UR�M�蟔���Kj h@�j�p�����E��}� t�EP�N�  ��P�MQ�M������E���E�    �U�R�M��t���E���]� ���������������������������������������������U��Q�M��M���k����tC�M��[l����u�}t�}u�EP�M��M�����} u��MQ��y����P�M��s���E���]� ���������������������������������U����M��M��`����uj�M��k����u^j h@�j�o�����E��}� t�EP�M��n���E���E�    �M�M�}� t �U�����E��M��U���E��M��U�T��E���]� ����������������������������������������U����M��M�������t3�M�j����u'�M�ۈ���E��E�%�   �M��Q�� ���ЋE��P�E���]� ������������������������������U��Q�M��E��M��U��E�B�M��A    �U��B    �E��@    ��]� ��������������������U��Q�M��E��x t7�M��U��B�A�M��y t"�U��B�M���Q�E��HQ�U��B�Ѓ��ɋ�]����������������������U���ٮ����t�E������M�����]������������������������U����M��} t_j h@�j�m�����E��}� t�EP�M��R�M��k���E���E�    �E��M��U��: u�E��H�� ������U��J��E��H�� ������U��J��]� ���������������������������������������U���  �M��^����k����E��M�<`���������}���  uj�M������E�8  �B�}���  u�EPj�MQ�Е�����E�  ��}���  u�UR�M�k���E��  �E�% �  �{  �M��� �  t5�U���   ��   uǅt���   �
ǅt���    ��t����������-�M��� `  uǅ����   �
ǅ����    ������������������ t�E�%   �E���M���   �M��}� tL�U��� �  t0�E�%   =   uǅ����   �
ǅ����    �������M���E�    �}� ��  �U��� �  t3�E�%   =   uǅ����   �
ǅ����    �������������$�U��� `  u	�E�   ��E�    �EЉ����������� t�M���   �M���U���   �Uȃ}� ��   �E�% �  t2�M���   ��   uǅ����   �
ǅ����    �������U���E�    �}� ��  �E�% �  t2�M���   ��   uǅ����   �
ǅ����    �������U���E�    �}� �q  �E�% @  tV�%\����t5������t,��p���Q�a����Pj ��`���R�������P�M��X���������P�la����P�M��r���M��� �  t5�U���   ��   uǅ����   �
ǅ����    �������������$�M��� `  u	�E�   ��E�    �U������������� t�E�%   �E���M���   �M��}� �O  �U��� �  t0�E�%   =   uǅ����   �
ǅ����    �������M���E�    �}� �  ������R�uh����P������Pj{�����Q�M�e�����ڀ��P�M��{���������R聫�����o����u4h����p���P������Qj,������R�}�����������P�M��/���h���M�苚��������P�t}�����SZ����tU�O}����tL�n����uC�M�Q��`���Rj ��P���P������Qj ��P���R�
��������~��������P�M��V���-
  ������臅���������|����������q����������f����������[����E�% �  t5�M���   ��   uǅ����   �
ǅ����    �������������#�E�% `  u	�E�   ��E�    �M������������� t�U���   �U���E�%   �E��}� ��  �M��� �  t5�U���   ��   uǅ����   �
ǅ����    �������������$�M��� `  u	�E�   ��E�    �U������������� te�E�%   =   uV������Q�t����P�������[U����@���R�t����P�������@U���� ���P�ot����P�������%U���   �M��� �  t,�U���   ��   u	�E�   ��E�    �E���x����-�M��� `  uǅ����   �
ǅ����    ��������x�����x��� t*�E�%   =   u��0���Q��s����P�������T��������R�s����P�������nT���E�% �  t5�M���   ��   uǅ����   �
ǅ����    ��������x����,�E�% `  uǅp���   �
ǅp���    ��p�����x�����x��� �  �U��� �  t3�E�%   =   uǅh���   �
ǅh���    ��h�����`����-�U��� `  uǅp���   �
ǅp���    ��p�����`�����`��� tS�M��� �  t5�U���   ��   uǅh���   �
ǅh���    ��h�����X����
ǅX���   ��X��� uA�w�����t�� ���Q�َ����P�������S�����@���R輎����P��������l���'V����tO�#y����t,�E�P�����Q������R�y�������
|��P�M��R����� ���P��x����P�M��l����� ���Q��x����P�M��il���M�`����uA�M��`����u)��i����u �URj ������P������P�M��8�����MQ�M��1R���E�    ����������������� tNj ������R舁����Ph��������P�f����P�M������ui����t�M�Q�M�Nb���E�  �ej h@�j�!c������`�����`��� t��`����x�����P����
ǅP���    ��P����U��E�P��0���Q������P�������cQ���U��� �  t3�E�%   =   uǅX���   �
ǅX���    ��X�����P����-�U��� `  uǅH���   �
ǅH���    ��H�����P�����P��� t�M���   ��@�����U���   ��@�����@��� ��  �E�% �  t5�M���   ��   uǅH���   �
ǅH���    ��H�����@����,�E�% `  uǅ8���   �
ǅ8���    ��8�����@�����@��� ��   �U���   ��   ��   j,������P������Q������Rj,������P������Q������Rj,��x���P������Qh����h���R��c�������w�����$y�����w�����y�����w��P�M�谡����   �E�% �  t5�M���   ��   uǅ0���   �
ǅ0���    ��0�����(����,�E�% `  uǅ8���   �
ǅ8���    ��8�����(�����(��� tG�U���   ��   u6j,��X���P������Qh���H���R�c��������v��P�M������h��M��L���h����8���P������胅��P�M��à��j)��(���Q�����R��f����Pj(�����P�׃�������lv��P�M�艠���M��� �  t5�U���   ��   uǅ0���   �
ǅ0���    ��0�����(����-�M��� `  uǅ ���   �
ǅ ���    �� �����(�����(��� ��   �E�% �  t5�M���   ��   uǅ���   �
ǅ���    �����������,�E�% `  uǅ ���   �
ǅ ���    �� ������������� tQ�U��� �  t3�E�%   =   uǅ���   �
ǅ���    �����������
ǅ���   ����� u������R�M��;����������t������P��^����P�M������������Q�^����P�M���f���Z����t������R������P�M��ߞ���������P������P�M��f��������Q�N}����P�M��f���q����t!�}� t�U�R�M��L��������P�M��L����  �MQ�M��r����U��� �  u,�E�% |  = h  u�M�Q�UR�_�����E�-  �  �E�% �  u.�M��� |  �� p  u�U�R�EP�O�����E��  ��  �M��� �  u]�U��� |  �� `  uLh���EP������Q��X����P������Rj{������P�M��s�����u�����_����E�  �g  �M��� �  u.�U��� |  �� |  u�E�P�MQ��V�����E�T  �.  �U��� �  t3�E�%   =   uǅ���   �
ǅ���    �����������-�U��� `  uǅ ���   �
ǅ ���    �� ������������� t�M���   ��������U���   ������������ td�E�% �  t5�M���   ��   uǅ ���   �
ǅ ���    �� ����������
ǅ����    ������ th,��M��ύ���-  �E�% �  t5�M���   ��   uǅ����   �
ǅ����    �������������,�E�% `  uǅl���   �
ǅl���    ��l��������������� t�U���   ��,�����E�%   ��,�����,��� te�M��� �  t5�U���   ��   uǅ����   �
ǅ����    ��������d����
ǅd���    ��d��� thT��M��Ό���,  �M��� �  t5�U���   ��   uǅ����   �
ǅ����    �������������-�M��� `  uǅ���   �
ǅ���    ����������������� t�E�%   ��\�����M���   ��\�����\��� t`�U��� �  t3�E�%   =   uǅ����   �
ǅ����    ��������$����
ǅ$���    ��$��� th���M��͋���.�U��� �  u#�E�% |  = x  u�M�Q�M�X���E�!	  �U��� �  t3�E�%   =   uǅ����   �
ǅ����    �������������-�U��� `  uǅT���   �
ǅT���    ��T��������������� t�M���   ��������U���   ������������ ��   �E�% �  t5�M���   ��   uǅ����   �
ǅ����    ��������L����
ǅL���    ��L��� uR�E�% �  t5�M���   ��   uǅ����   �
ǅ����    ������������
ǅ���    ����� t#�E�Ph����x���Q��Z����P�M���F����U�R��h���P�,V����P�M��F���M��� �  t5�U���   ��   uǅ����   �
ǅ����    �������������-�M��� `  uǅD���   �
ǅD���    ��D��������������� �#  �c�����   �E�% �  t5�M���   ��   uǅ���   �
ǅ���    �������<����,�E�% `  uǅ����   �
ǅ����    ��������<�����<��� tr�U��� �  t3�E�%   =   uǅ����   �
ǅ����    ������������
ǅ���   ����� t!�U�Rh̼��X���P�eY����P�M��JE���M��� �  t�U���   ��   ��  �E�% �  t2�M���   ��   uǅ|���   �
ǅ|���    ��|����U��)�E�% `  uǅ4���   �
ǅ4���    ��4����M�}� t�U���   ��������E�%   ������������ �c  �M��� �  t)�U���   ��   u	�E�   ��E�    �E�E��!�M��� `  u	�E�   ��E�    �U�U܃}� t�E�%   =   ��   �M��� �  t)�U���   ��   u	�E�   ��E�    �EԉE��!�M��� `  u	�E�   ��E�    �ỦUă}� t�E�%   =   tj�M��� �  t)�U���   ��   u	�E�   ��E�    �E��E��!�M��� `  u	�E�   ��E�    �U��U��}� t0�E�%   =   u!�M�Qhؼ��H���R�KW����P�M��0C���q������	  �E�% �  t)�M���   ��   u	�E�   ��E�    �U��U�� �E�% `  u	�E�   ��E�    �M��M��}� ��   �U��� �  t(�E�%�   ��@u	�E�   ��E�    �M���|����*�U���   ��   u	�E�   ��E�    �E���|�����|��� t&�M�Qh���8���R�ZV����P�M��?B���   �E�% �  t5�M���   ��   uǅt���   �
ǅt���    ��t�����d����,�E�% `  uǅl���   �
ǅl���    ��l�����d�����d��� ��   �U��� �  t3�E�%�   =�   uǅ\���   �
ǅ\���    ��\�����L����3�U���   ��   uǅT���   �
ǅT���    ��T�����L�����L��� t&�M�Qh���(���R�BU����P�M��'A���  �E�% �  t5�M���   ��   uǅD���   �
ǅD���    ��D�����4����,�E�% `  uǅ<���   �
ǅ<���    ��<�����4�����4��� ��   �U��� �  t.�E�%�   uǅ,���   �
ǅ,���    ��,���������-�U���   uǅ$���   �
ǅ$���    ��$������������� t!�M�Qh ������R�5T����P�M��@���E�% �  t5�M���   ��   uǅ���   �
ǅ���    �����������,�E�% `  uǅ���   �
ǅ���    ��������������� t�U���   ��������E�%   ������������ t*�W����u!�M�Qh������R�oS����P�M��T?���E�%   t!�M�Qh�������R�DS����P�M��)?���E�P�M�O���E��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�M�jPh`��M��y���`���]������������������U��Q�4�%�   u	�E�   ��E�    �E���]����������U��Q�4���u	�E�   ��E�    �E���]������������U��Q�4���u	�E�   ��E�    �E���]������������U��Q�4�% �  u	�E�   ��E�    �E���]����������U��Q�4�%   u	�E�   ��E�    �E���]����������U��Q�4���u	�E�   ��E�    �E���]������������U��Q�4���u	�E�   ��E�    �E���]������������U��Q�4�%   u	�E�   ��E�    �E���]����������U��4�%   ]������������������U��4�%   ]������������������U����M��E��8 tj�M��]���  �} ��   �} ��   �M�M��}� t�}�t�u�U��B% ������M��A�   j h@�j��F�����E�}� t�U�P�M��y���E���E�    �M��U���E��8 u�M��Q�� ������E��P�[j h@�j�F�����E�}� t�MQ�UR�M���j���E���E�    �E��M��U��: u�E��H�� ������U��J��E��H�� ������U��J��]� �������������������������������������������������������������������������������������������U��Q�4�%   u	�E�   ��E�    �E���]����������U��Q�4�%   u	�E�   ��E�    �E���]����������U��Q�4���`��`t	�E�   ��E�    �E���]�������������������������U��Q�4�%   u	�E�   ��E�    �E���]����������U��4�%    ]������������������U��Q�4���u	�E�   ��E�    �E���]������������U���,�E�   �M��b���M��^�����  �$����@��   �$����Z��   �}� t	�E�    �
j,�M��T���$������   �$����0�M�x3�}�	-�$����$��E�P�M�Q���5��P�M�蚄���k�$��U�M��ia��P�E�P��Z�����$�+M��~����4����u�U�R����1���E�P�M��B����$�;M�u
j�M���Y���j�M��2����������U�R�M�B���E��]�������������������������������������������������������������������������������������������U��� �$���M��}�XtD�}�Zt�`�$����$���Y����t	�E�Pl��E��E�P�M�Z���E��   �$����$�h̻�M�6���E��   �U�R�V�����M��\������   �$���M��}� t�}�@t`�}�Zt�v�U�R�M�lA���E�   �$����$��NY����t	�E���E��M�Q�U�R�M��bg��P�M�%A���E�>�$����$��M�Q�M�A���E� j�M�o���E���U�R�M��@���E��]�����������������������������������������������������������������������������������������������U���   �$�����~  �h:���E��}� }�E�    �}� u>j]�U�Rj�E�Pj[�M��#q�����.P�����W��P�MQ�B�����E��  �   �M��e^���M��i����th���M���r���M��z<����tZ�U��U��E����E��}� tE�$����t8j]��x���Pj �M�Q�l����Pj[�U�R�Td��������V��P�M�����뚋M�<����ua�M�Di����t�E�P�M�Q�M�2X��P�M���.���:�U�R��h���Pj)�M�Q�URj(�E�P��c�������V������W��P�M��.���M�Q�U�R��V�����M���O���E�P�M��>���E�   �   �M�<����uPj]�M�Qj�U�Rh ��E�P�MQj(�U�R�qc��������d�����N������U��P�EP�0A�����E�<�:j]�M�Qj��p���Rj[��`����^o�����iN�����U��P�EP��@�����E��]������������������������������������������������������������������������������������������������������������������������������������������������U���j �[����P�M��#{���$����tl�$���E��$����$��U��U��}�0t�}�2t�}�5t(�5h̻�M��?p���&�E�P��;����P�M��~���j�M�]k���E�(�
j�M��|��h(��M���o���M�Q�M�=���E��]������������������������������������������������������U���t�$�����k  �$���E��$����$��E� �E������M���Z���U��U�E��C�E�}��   �M���x��$�L�h���M��!a���?  hȽ�M��a���-  hн�M���`���  hԽ�M���`���	  hܽ�M���`����  hD��M���`��h��M���n����  �E����E���  �$���U��E��E�$����$��U�U�}�Y�8  �E������$����E������(  h��M��K`���  h���M��9`���  h���M��'`����   h��M��`����   h��M��`����   h ��M���_���   h,��M���_���   h8��M���_���   �$����$��E�P�1����P�M��\*���M���7����t�M�Q�M��:���E�~  �R�UR�E�P�B=����PhD��MQ�*>�����E�R  �$����$�j�M��Q���hL��M��0_���Qh̻�M��!_���B�$����$��M�Q��0����P�M��)���M��O7����t�U�R�M�:���E��  �}����   �E��E��M���C�M��}���   �U���8��$�(��M�QhL��U�R�]=����P�M��B)���e�E�PhX��M�Q�==����P�M��")���E�U��U�E��E�E�}�w/�M���`��$�X��E�PhL��M�Q��<����P�M���(���M�u6����u�URj �E�P��]����P�M��z���M�Q�M�$9���E��   ��   �M��nW���UR�M��9���}��uF�M���I���E�P�M�Q�U�R�pa�����M��b����uh���M��k���E�P�M�8���E�}�M��5����tA�M���t$hd��M��b]���U���thl��M��gk����E���th`��M��6]���M�Q�U�R�EP��5�����E���MQj�UR�\b�����E��]Ë��0�B�T�f���x������-�   










	�I ������*�<�N�����`�r���� 	
��������)� �I �)�     ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP��a�����E]�����������U����$�����0  �$����A�E��$����$��}���   j�M��_c����'������   �U�����U��}���   �E���|��$�X�j��R����P�M���Y���   j��R����P�M��Y���|j�R����P�M��Y���gj�R����P�M��~Y���Rj�R����P�M��iY���=j�vR����P�M��TY���(j�aR����P�M��?Y���j�LR����P�M��*Y���U�R�M�R4���E� �j�M�hb���E��j�M�Wb���E��]Ðy��������������"� ���������������������������������������������������������������������������������������������������U���0  �M���Q���E� �$�����5  �   k� �$����$u8�EP�M�Q�UR�E�P��*�����M��Z0����u�M�Q�M�$3���E�  �$����A|	�E�A   ��E�   �$��+UԉU��M��FQ���M��>Q���E�   �E��E��}�t�}�tw�}���   �#  �t%����tZ��b����tQ�M���/����u2j	�tP����P������Qj �U�R�M���I�����X��P�M���!���j	�BP����P�M�� W����   �%����tQ�M��d/����u2j�P����P������Pj �M�Q�M��qI�����GX��P�M��!���j��O����P�M���V���f�$����tT�M��/����u5j
�O����P��(���Rj ��x���P�M��I������W��P�M��/!���j
�O����P�M��bV����E�    �}� ��   �$����$��   k� �$����$u8�EP�M�Q�UR�E�P�)�����M��c.����u�M�Q�M�-1���E�  �$����A|	�E�A   ��E�   �$��+UЉU��}� �����$����t�$����$��}��|  �EP�M��9n���M�Q�U�R�M��I��P�M��( ���M���-����u,�E�P��h���Qj �����R�M���G�����HI��P�M������M��-����u,�E�P��X���Qj ������R�M��G�����I��P�M�����E����  �} tj�M�?^���E�  �M���tw�E�PhT���H���Q�3����P�M��i���$����t,�M�Q�����R��8���P�D�������H��P�M��2����M�Qj�U�R�Y����P�M�����!�$����t�U�R�LD����P�M���8���$����uj�M���n���3�$���E̋$����$��}�@tj�M�R]���E�  ��!����tR�U����Uȃ}�t�?�} tj�M� ]���E�q  �E�P�M�Q��p���R�+'�������G��P�M��N���#�E�����u��`���Q��&����P�M��8���U���t!�E�Ph̾��P���Q�2����P�M�� ���U���t!�E�Phؾ��@���Q��1����P�M������} ��   �M�g+������   �M�Y����u�M�K+����t:�M��W����t�UR�M������EPj ��0���Q�R����P�M��fo���@�UR�� ���Pj �����Q�URj �� ���P�yR�������E�����F��P�M��$o���*�M��*����u�MQj ������R�?R����P�M���n���M���+���E���t�M��uR���M�Q�M�W-���E��   �j�M�j[���E�   �   �} ux�M�N*����ul�M�X����u�M�6*����t�URj�EP�W�����E�u�9�MQ�URj ������P�MQj������R��V�������D�����E���E�:�8�} u%�M��)����u�EPj�MQ�V�����E��j�M�Z���E��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E��Qj �M���H��P�E�P�M���H��P�MQ�\<�����E��]�������������������������U��� �EP�M���)���$���U��}� t�}�?tq�}�Xt��   �E�Pj�MQ�9T�����E��   �$����$��M��!'����th̻�M�fg���E�   ��E�PhX��MQ�a-�����E�w�$����$��E��Qj �M��H��P�E�P�M�Q�U�R�n;����P�M�����E�P�MQ�^A�����E�$�U�R�M�g)���E��E�P�MQ�8A�����E��]����������������������������������������������������������������������������U���h�C+����tH�4�%�����4�j �M�Q�������4���    �4��E�P�M�(���E��  ��  �$����?��  �$����$��   k� �$����?uS�   �� �$����?u=�U�R�u!�����$����t�$����$���E�P�M�)(���E�9  �M�Q��G�����M��Z���E��M��� ���E��M��$����u�U�R�M��'���E��  �$������   �$����@��   �M�Q�<�����M���$������   �8���tn�8� �E�P�M�Q�M��R@��P�M������$����@t>�M�Q�1<����P�M������U�R�E�PhT��M�Q�M��nM�����@��P�M�����)�U�R�E�PhT��M�Q�M��CM������?��P�M�����}� t�M��t&���}� t�M��-���M��$����u�M��>&����t�U�R�M�&���E��   �   �$����t�$����@ut�$����t�$����$��-����t:�}� u4�M��A����u(�M��D��P�M�Q�3�����U�R�M�B&���E�U��E�P�MQ�3�����E�>�j�M�AT���E�-�+�$����tj�M�#T���E��j�M�T���E��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   V�E�    �$����Qu�E����$����$��$����uj�M��R���E�W  �R  �$����0��   �$����9��   �}� tG�$�� ��/��EЉUԋ$����$��U�R�E�P�M��V��P�M�Q�U�R��'�����E��4�$�� ��/��EȉŰ$����$��U�R�E�P�M���U���E��M��M�U�R�M�$���E�  �  �E�    �E�    �$����@��   �$����uj�M��Q���E�P  �W�$����A|7�$����P*�E؋Uܱ�Vd���ȋ�$����A���M؉u��j�M�Q���E��   �$����$��e����$���U�$����$��}�@tj�M�JQ���E�   �M��tX�}� t&�U�R�E�P�M��T��P�M�Q�U�R�&�����E���E�P�M�Q�M��T���E�U�U�E�P�M��"���E�V�T�}� t&�M�Q�U�R�M��dT��P�E�P�M�Q�*&�����E���U�R�E�P�M��>T���E��M��M��U�R�M�j"���E^��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�$����tw�$����_ui�$��Q��t[�$��H��_uM�$����$��$����$��$����A�U��$����$��}�vj�M�UO���E��M�?���E��]�������������������������������������������U��j�EP�GM�����E]�����������U���8��S����t��'����u	�E�   ��E�    �E��E�M���>���$���U�$����$��M��M��}�Y��   �U��� �$� �$����$�hy��M��]���E�   h���M���D���kh���M���D���\h���M���D���Mh���M���D���>h���M��D���/��R���E�U�R�,����Phľ�E�P�a#����P�M��F���M��>���}� t�M�Q�M��,���U�R��^����P�M��a���E�P�M����E��]� DSb�q�� ����������������������������������������������������������������������������������������������������������������������U��EP�!�����E]�������������U����M���<���$������   �$���E��M���0�M��}�wH�U��$�$h,��M���B���>h4��M���B���/�-h<��M���B���hD��M��B���j�M�L���E�~�$���M�$����$��E�E��M���1�M��}�w/�U���L�$�D�M�QhL��U�R�!!����P�M�����E�P�M�v���E��j�M�K���E��]Ë�SSbbqs����    ���������������������������������������������������������������������������������������������U���0�M��!;���$����$��$���U��}�At�}�BtU�}�C��   �   �} u,�E����&u	�E� ���M����*u	�M���$����$��  �} tj�M�`J���E�  �E� j>�M��#���$����$��p  �U����$����$��U  �   k� �$����t�   �� �$����uj�M��I���E�$  �} tj�M��I���E�  �   k� �$����0���   �� �$���LЉM��$����$��}�v/j,�M��8"���E�3�QP�M���L��P�U�R�M��4��P�M��
��j>�E�P�M��r2��P�M��
���$����$u�$����$��j^�M�Q�M��>2��P�M��b
���$����t�$����$��
j�M��DZ���M��)���U�R�M����E��M��8���E��]���������������������������������������������������������������������������������������������������������������������������������������������������������������U���,j h@�j�������E��}� t�M��'8���E���E�    �E��E�M�Q�U�R�	�����EP�M�Qj �U�R�E�P����������0�����Q2��P�M������M�Q�M�i���E��]���������������������������������������������������U����   �$����u�URj�EP�(C�����E�/  �$����6|�$����9~ �$����_tj�M��F���E��  �$����6�U��$����$��}�)u[�$����t2�$����=�M��$����$��}�|�}�~�E�������EPj�MQ�rB�����E�y  ��}� |�}�~�E������}��uj�M�MF���E�L  �M��u6���UR�M��
���E����  �M�QhT���X���R�|����P�M��a���$����t;�U�R��H���P�M�Q�,����Pj ��h���R�c<�������t0��P�M������E�Pj�M�Q�A����P�M������$����t1�$����@u�$����$��j�M�nE���E�m  ��M�Qj�UR�JA�����E�Q  ��Y����t��(���P�QB����P�M������M�Q�:B����P�M��Z ���U���tY�	����t8�E�P�M�Q�U�R�����Pj ��8���P�o;�������/��P�M��(�����x���Q������P�M������G	����t&�U�R�E�P�M�Q�K,�������9/��P�M�������U�R�-,����P�M�����M�d����u(j)�E�P�M�Qj(�U�R��:�������r-��P�M����j h@�j�������E�}� t�M��O4���E���E�    �E�E��M�Q�U�R��4����j)�E�P��p���Q�Z����Pj(��`���R�b:��������,��P�M��W���cX����t�E���t�M�Q�M���V���>����t��P���R�����P�M���V�����@���P�h����P�M����������t��0���Q��8����P�M��V����� ���R�8����P�M��s���}� t�E�P�M��v���j�M�C���E��M�Q�M�����E��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�@�����E]�����������U��Q�M��M������t2���E���U���
�P�ҋ�]���������������������U����M��E��xu�   k������E���E� �E���]�����������������U��Q�M��E��@��]����������������U����M��E��x t�M��I�9���E���E� �E���]��������������������U����M��E��H�U���J�P�҈E��E���u�M��Q�E���H�B�ЈE��E���]�����������������������������U����M��E��x t�M��Q�E��H�T��U���E� �E���]���������������U���j'�EPj �M�Q�^>����Pj`�U�R�6�������7)���E��]��������������������������U����M��E������E�} t�MQ�U���Ѓ���   ��   �} w�E   �M��Q;U��   �}   v3��   jh@�h  �;�����E�}� t�M�����E���E�    �E��E��}� tA�M��y t�U��B�M���U��E��B��M��U��Q�E��M��H�   +U�E��P�3��!��M��Q+U�E��P�M��Q�E��H�D
��]� ������������������������������������������������������������������������U����$����u3���   ��   �$����0|8�$����9*�$����/�M��$����$��E��   �   �E�    �$����@tY�$����u3��o�7�$����A|$�$����P�U����$���T
��U������6�$����$�뚋$���U��$����$��}�@t�����E���]���������������������������������������������������������������������U���  �M��~-���M��v-���E�    �E�    �$���M��$����$��E��EЃ}�_��  �M����*�$��*�$����$�j�M��<���E��  �M��-���M����   ��<���R�����Pj<��l���P�53����P�M���O���M������ȃ�>u
j �M����j>�M�����} t�U��$����u�U�R�M�)���E�>  �$����$��$��M�j j ��,���R��7����P�M��s����E��$��M������u4�   k���$����1u�U�Rj~��\���P�k2����P�M��+����M���
����u�M�Q�M��O���U�R�M����E�  �G  �   k���$��
��P�Q�M�� 2���   �E�   �   k���$����4�P�M���1����  �$���U��$����$��M��Mԃ}�_��  �U���T+�$� +�$����$�j�M��:���E��  �   k���$�����P�M��p1���_  �   k���$�����R�M��I���E�  �1  �   k���$��
���Q�M���I���M�����U�R�M�;���E�P  ��  jhd��E�P��������M��1���M�Q�M����E�  �   k���$����ĲP�M�YI���E��  �   k���$����ĲR�M��0��j j �����P�q����P�M������M������u�M���(����tj�M�9���E�  �M�Q�UR�M��1$���E�s  �  �  �   k���$��
��ĲQ�M���/���   k� �$����uj�EP�M�����E�  �   k� �$����0�M�x�}�rj�M��8���E��  �U���X�P�M��/���$���U��$����$��M��M�U��0�U�}��;  �E��$��+j �M�Q�e������U�R�EP�M�Q��L���Rj �����P�M��!�����#�����#���E�S  �  �M�Q�U�R�M���"��j,��|���P������Q��������Y!��P�M��vK��j,��t���R��d���P���������1!��P�M��NK��j,��T���Q��D���R��������	!��P�M��&K��j)��4���Pj ��$���Q��5�������� ��P�M���J��j'�UR�M��� ���E�  �;�E�P�MQ�M��*"���E�l  �!�$����$�j�M�[7���E�I  ��  �   k���$��
��ĲQ�M���-����  �$���E��$����$��U��U؃}� t�}�0t!�N�$����$�j�M��6���E��  j h���M�Q�a������M��.���U�R�M����E�  j�M�6���E�  �,  �$���M��$����$��E��E�M��A�M�}�	��   �U����+�$��+�   k���$����(�R�M�E���E�  �   k���$��
��(�Q�M��YE���$����?u7�����Q�� ����P�M��4I���$����@u�$����$�������R�q'����P�M���H��h���M��Y:���E�P�M�g���E��j�M�}5���E�n�j�M�l5���E�]�j�M�[5���E�L�}� t
�M�����-�M��=����u!�M�Qh��������R�
����P�M��v����E�P�M�����E��]ÍI �"�"
$8$1$_$B* �$�$�$%�(�%R%�%/&4&Y()1* 	

'O'(((X)�)        ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�E�4p�E�P�MQ�UR�EP��-�����E��]�����������������������U��Q�E��Q�E�P�MQ�UR�EP�-�����E��]�����������������������U���<�M��!���$���M��}�B��  �U����1�$��1�MQj�UR�,�����E�s  h`��M��1'���M������u
j �M�����EP�M��C���$����$��E����U�R�M�� ��P�E�P�MQ�2�����E�	  �   �� �$����$tC�   �� �$����u�URj�EP��+�����E��  �j�M��/���E�  �$����$��$���E��}�T�i  �M���2�$��1�$����$��MQ�UR�!�����E�U  �$����$�j�MQ�UR�@�����E�.  �$����$��E��Qj �M��n��P�M�Q�UR�E�P������P�MQ������E��   ��   h`��M��%���M�������u
j �M������UR�M�� ���$����$��E���M�Q�M�����P�U�R�EP������E�|�$����$�j�M�.���E�^�I�$����$�hl��M�=���E�;�&�EPj�MQ�E*�����E�"j�M�>.���E��UR�EP������E��]ÍI �.x/1//n1 �H10,0S0�0�01%1_1 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����$�����  �} t]�$����XuO�$����$��M�%�����th̻�M�j;���E��   ��URhX��EP�e�����E��   �$����Yu%�$����$��MQ�UR�I������E�   �EP�M�Q�  �����M������t �U�Rh��E�P�� ����P�M�������*�M�e)����t�M�Qh��U�R�� ����P�M������E�P�M�"����E���MQj�UR�('�����E��]�����������������������������������������������������������������������������������U����$������   �$����6|�$����9~�$����_un�UR�M���9���M������u$�M�w�����u�M�'����u�EP�M��=���M�S�����u�MQ�M��=���U�R�EP�������E�   �Nj �MQ�UR�EP�M�Q�������U���*u	�E�   ��E�    �M�Q�U�R�EP�(;�����E�m�kj�M���)���MQ�M��.���M������u�UR�M��=���M������u"�M������u
j �M�����EP�M���<���M�Q�M�K����E��]�����������������������������������������������������������������������������������������������������U��EP�MQ�UR�EP�%�����E]�����������������U����$�����  �$����_�  �$����$��$����A�E��$����$��}���   �M������������   h���M��-��j�
����P�M��-���}� tk�U��҃�#U��U�E�E��}�t�}�t�h���M���,���h���M��,���j�M��'���E�U�M���#M��M�th���M��,���j)�M���
���U�R�M�����E��j�M�'���E���M�����E��]�����������������������������������������������������������������������������������������������U��$����@u"�$����$��EP�M�����E���MQ�UR��������E]��������������������������U����   �M������E� �M��x������  �$������  �$����@��  �8���t�9���u�E�P�M�G����E�-  �M��]�����uH�M�QhT��U�R������P�M������E���t"�M�Qj[��d���R�����P�M��s����E� �$����?�  �$����$��$���M��U���$�U��}�-��  �E����=�$�t=�   �� �$����_um�   ��$����?uX�$����$��E�P�M�Qj j ��4���R����������P�M������$����@u�$����$��F�E�P�M�Qj'��T���R�E�P������Pj`�����Q��������:�������P�M��W�����  �$����$��E�P�M�Qj j��D���R� �������p��P�M������  j@h$��M��&���E�Ph����t���Q�������P�M���������:�����u�U�R���k����l  �$����$��M�Q��$���Rj]�E�Pj j�M�Q���������^��������P�M��{����E��  �M��E���$����$�j j�E�P������M������uE�M��������u+�M�Q�U�RhT��E�P�M��������b��P�M��
�����M�Q�M�������
j�M�����M��I����u�$����@�w����M��+����u<j]�M�Q�U�Rj[��|���P���������w��P�M������$����$��
j�M��0���*�U�R��l���P��\���Q����������P�M��T����.�U�R��L���Pj j��<���Q��������|��P�M��$���� ����$���E�}� t�}�@tW�W�M�������tj�M�����;�M�Q��,���RhT������Pj������m"�����s�������P�M�������
j�M��U���M�Q�M�����E��]Ë��:�:�9D;�;�< ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���@�M�����j j�E�P�E����P�M�������M��6����uN�$����tA�$����@t4�U�R�E�PhT��M�Q�U�R���������C������
��P�M������$����@u�$����$��b�$����tj�M������J�M��������tj�M������2�U�R�E�PhT��M�Qj�M�������������[
��P�M������U�R�M�s����E��]�����������������������������������������������������������������������������U����$����uj�M�+���E�T�R�$����?u3�$����$�j �U�R�:����Pj-�EP�~�����E��j �MQ������E��]����������������������������������������U��EP��������E]�������������U��Q�M��M��w�����t�E��EP�MQ�U���M���	�B�Ћ�]� �������������������������U����M��M��%�����uX�} u*�M���(�����Ej h@��EP��������E��M��M�} t �U�E�L�Q�UR�M��{"���E�E��  ��} t�M� �E��]� ����������������������������������������������U��Q�M��E��xujh���MQ�UR�Q*������E��]� ��������������U��Q�M��E;Es�M�U��B��M���M�E��]� ��������������������U����M��E��x t�MQ�UR�E��H�!���E���M�M��E���]� �����������������������U����M��EP�MQ�U��B�M���I�B�ЉE��M�;Ms�UR�E�P�M��Q�E���H�B�����E���]� �������������������������U��Q�M��E��HQ�U��BP�MQ�UR�)������]� ���������������������U��� �EP�M��J+���$���U��$����$��}�@u�$���U��$����$��}�_tj�M����E�   �$����$�j �U�R������j �E�P������$����t�$����@t�$����$��ա$����u�$����$�j�M�*���E��$����$��M�Q�M������E��]�������������������������������������������������������������������������������U��Q�E+E�E��M;M�~�U��U�EP�MQ�UR�'  ���EE��]������������������������U��   k� �$��
��?uR�   �� �$��
��$uj�MQ��������E�;�$�$����$�j j �EP�������E��j j�MQ������E]������������������������������������������������U���|���3ŉE��E��M���	���9��M��J������  �$������  �$����@��  �E� �M��t�E� ��E��$����0�E�x6�}�	0�$����$��U�R�E�P� ��E���P�M��`,���<  �$��MčM��,	���E� �$����$uT�$��Q��$uE�$��H��Wu�E��$����$��"�$��H��Vu�$����$�������$����Xu!�$����$�h̻�M��
���,  �$����$u?�   �� �$����$t)�$����$��E�P�:�����P�M��v�����   �$����?��   �E�P��������)�����tkj�M�Q�M������U�R�4#����P�<����EЃ}� t�E�P�M��Y���.h���M�Q�U�RhԻ�E�P�����������P�M�������.h���M�Q�U�RhԻ�E�P����������j��P�M�������M����P�M�Q�� ����P�M������$�+Uă�~� ��������u�E�P� ������M��������u3�M��t
j,�M�������U�R�M��4*���E��thPl�M�����0����9� �M�Q�M�����E�M�3��V�����]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���  ���3ŉE��$���M��$����$��E���l�����l���T��  ��l�����LN�$�$N�EP�F������E��  �$����@u$�$����$�h��M�$���E�  �3�����Q�'�����P�URh����D����k$���������E�t  �EP��������E�`  ��T���Q��������\���R��������T����8�������   ��\����%�������   jd�   �� �L�Q��T��������uj�M����E��  �   �� �   k� �T��T��   k� �T���-u%�   ��   �� �T��T��   ���D�.��   �� �D�.��\���R�EPje������Q�U�R�������U#�����)����������E�W  �j�M�����E�C  ��d���P�������������tMj�M�Q��d��������U�R�����P�<�����p�����p��� t��p���P�M��"���E��  �M���Du5h���UR��d���PhԻ��,���Q���������J���E�  �3h���UR��d���Ph�������Q�~�����������E�m  �h  j j ��L���R����������P��������L���Q�M�����E�/  j{��x����{���U���t�����t���H|3��t���J~�(��<���P������P��x�����%��j,��x��������M��M��U���F�U��}�wu�E��$��N��4���Q������P��x����%��j,��x����;�����$���R�������P��x����c%��j,��x������������P�������P��x����;%��j}�MQ��x��������E�<�:�M�����E�-�+�$����$�j�M����E�j�M����E�M�3��;�����]Ë��M'J;J�J�K�J�L�L�MN 																																																																						�I MWM�MMWM����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   �   k� �$��
��?u�   �� �$��
��$tj�M�f���E�|  �$����$����U���E�� ��M�M�������h���������<��������U�����h�������<���� ��M��'����M������E� �$����?u,�$����$��U�Rj�E�P�]�����P�M������jj�M�Q�U
����P�M�������M�������t�8��U���uj�E�P�f�����Pj<�M�Q������P�M��!���M������Ѓ�>u
j �M��J���j>�M��@����E��t�$����t�$����$��M���U����E� ��M�Q�M�����E��]������������������������������������������������������������������������������������������������������������������������U����E��Qj�M�����P�E�P�M��{���P�MQ��������E��]�������������������������U���(�$����tg�$����Zu'�$����$��M�����P�M�����E�^�0j)�UR�E�P�8�����Ph���M�Q��������������E�,�*j)�URj�E�Ph���M��������V����������E��]������������������������������������������U���x�E�    �$����_u�U��� @  �U��$����$��$����A�  �$����Z�  �$����A�E�$����$��U��� �  �U��E��t�M���    �M���U��������U��}���  �E�% �  t�M���������   �M��U��U���E�%�����E��M��M��U���U�t�}�t@�}�tq�   �E�% �  t�M���?�����@�M���U���������   �U�E�E��r�M��� �  t�U���?����ʀ   �U���E�%����   �E��M��M��;�U��� �  t�E�%?����E���M��������M܋U܉U���E���  �E��k  �E���E؃}���   �M��$�t\�U���������   �U��   �E�%����   �E��s�M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��MԋUԉUЋEЉE����E���  �E��  �  �$����$��  �E� �$����$��$���Ũ}�R�]  �E����\�$��\�U����d���� �  �U��D  �E�%�g�� �  �E��/  �M����d���� �  �M��  �U����d���� �  �U��  �E�%���� |  �E���  �$��Q��Pu�$����$��$����$��$���Eȃ}�Q��   �M��� ]�$�]�$����$�����  �$����$��$����0|C�$����95�$���$��D
ѣ$������E��M���   �M��E��-  ��E���  �7�$����$�����	  �E���  �E���  �E���  �E���  ��  �E���  �$����$���  �E��$����$��$����0|�$����5~$�$����t	�E���  ��E���  �E��z  �$����0�EċM��� �  �M��U��� �  t�E�%����   �E��M��M���U��������U��E��E��M���t�U���������   �U���E�%����   �E��Mă�t�U���    �U���E�%�����E��Mă��M�t�}�t@�}�tr�   �U��� �  t�E�%?�����@�E���M���������   �M��U��U��s�E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��;�M��� �  t�U���?����U���E�%�����E��M��M���E���  �E��  ��E���  �E��  �$����$���  �$����0��  �$����8��  �$���U��$����$��M�������M��U��U��E���0�E��}��?  �M��$�t]�U��� �  t�E�%����   �E��=�M��� �  t�U���������   �U��E��E���M��������M��U��U��E��E��M��M��U��� �  t�E�%?�����@�E���M���������   �M��U��U��  �E�% �  t�M���������   �M��;�U��� �  t�E�%����   �E��M��M���U��������U��E��E��M��M��U��U��E�% �  t�M���?����ɀ   �M���U���������   �U��E��E��  �M��� �  t�U���������   �U��;�E�% �  t�M���������   �M��U��U���E�%�����E��M��M��U��U��E��E��M��� �  t�U���?����U���E�%�����E��M��M��   �U��������� @  �U��l�E�%���� `  �E��Z�M���������    �M��F�U��������� h  �U��2�E�%���� p  �E�� �M��������� x  �M���E���  �E��H�C�$����9u�$����$��E���  ��$����t	�E���  ��E���  �E���]Ð�U�UJU�U8U�U!U�W{V�WV#VfV8VOV�WXY 																																																																					�fW�V�VMWuW ���Y~Z[�[�[�[�[�[\����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�$���M��}� t)�}�At�0�$����$�h��M����E�j�M�0����E�j�M�!����E��]������������������������������������U��EP�MQ�������E]���������U����EP�M�����h��M��w���M�Q�Z�����P�M�����j}�M������$����@u�$����$��U�R�M�I����E��]�����������������������������������U���@�EP�M������M��������b  �$�����Q  �E�P�M�Qj �U�R�E�P�'��������#���������P�M��@����M��I������  �$����@��   h��M��s���M���������   �$������   �$����@txj'�M�Q�U�R�"�����Pj`�E�P�������������P�M�����$����@u�$����$��M�������t�$����@th��M������Z����M��t�����t �$����u
j�M��S��j}�M�������$����@u�$����$��'�M��)�����t�U�Rj�E�P������P�M�������M�Q�M�i����E��]�������������������������������������������������������������������������������������������������������������������U���p���3ŉE��$����0�M�x5�}�	/�$����$��E�P�MQ�������E�N  �I  �M�������$����?utj �M�Q�F�����P�M������$���Eȋ$����$��}�@t7�$����$��$����t	�E�   ��E�   �U�R�M��J����  jhX��$�P��  ����u�E�X��$����$��7jhp��$�R�  ����u�E�p��$����$���E�    �}� ��   �M�Q�������������twj�U�R�M�������E�P������P�<����E؃}� t�M�Q�M������:h���M�����h���U�R�E�P�M�Q�U�R���������R���P�M�����:h���M������h���E�P�M�Q�U�R�E�P������������P�M��V���P�M��t0�$����@u"�M�����P�M��4����$����$��j@h$��M��.���P�M������U��t���Z�����u�E�P��苺���M�Q�M�U����E�M�3��!�����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��4�% @  ]������������������U��Q�M��E��@������]����������U��Q�M��E��@������]����������U����M��E��8 u	�E�   ��E�    �E���]�������������������������U����M��E��8	u	�E�   ��E�    �E���]�������������������������U��Q�M��E��@������]����������U��Q�M��E��@������]����������U��Q�M��E��@������]����������U����M��M��e�����u�E��H��	��t	�E�   ��E�    �E���]�����������������������U����M��M�������u�E��H��
��t	�E�   ��E�    �E���]�����������������������U��Q�M��E��@������]����������U����M��E��H������	�E�   ��E�    �E���]����������������U��Q�M��M��g�����t3���E���U���
��ҋ�]����������������������U��Q�M��E��@��]����������������U��Q�M��   ��]�����������������U����M��E��x t�M��I� ���E���E�    �E���]�����������������U��QV�M��E��x }.�M��Q�E���H��Ћ��M��Q�E���H�����M��q�U��B^��]�����������������������U��Q�M��E��@��]����������������U��j�h�d�    P���3�P�E�d�    �����uM���������E�    j ����"���j�������j����
���j���������E������} |�}}kE����   k����M�d�    Y��]�����������������������������������������������������U��Q�M��E��H��   �U��J��]��������������������U��Q�M��E��H�� @  �U��J��]��������������������U��Q�M��E��H��   �U��J��]��������������������U��Q�M��E��H��    �U��J��]��������������������U��Q�M��M�������u�E��H��   �U��J��]������������������������U��Q�M��E��H�� �  �U��J��]��������������������U��Q�M��E��H��   �U��J�E���]�����������������U��Q�M��E��@������]����������U��Q�E�    �	�E����E��M�;Ms�UU��EE���
�݋�]�����������������������������U��Q�E�    �	�E���E�M���t�E����E���E���]���������������U��} u3��G�E���Et.�M���t$�E��U�;�u�M���M�U���U�ǋE� �M�+�]���������������������������U��j�h�h�Ld�    P�ĜSVW���1E�3�P�E�d�    �} u3��   �E�    j�5������u3��oj�T������E�    �EP�MQ�@�������URj �EP�MQ�UR�M�������M������E�@������E������   �j�V�����ËE�M�d�    Y_^[��]����������������������������������������������������������U��j�h(�h�Ld�    P�ĜSVW���1E�3�P�E�d�    �} u3��   �E�    j�%������u3��pj�D������E�    �EP�MQ�@�������U R�EP�MQ�UR�EP�M�������M������E�@������E������   �j�E�����ËE�M�d�    Y_^[��]���������������������������������������������������������U��W�= ���   �}ww�U�����fn��p� ۹   #σ����+�3��of��ft�ft�f��#�uf��#���ǅ�EЃ������Sf��#���3�+�#�I#�[��ǅ�D�_���U��t93���   t�;�Dǅ�t G��   u�fn�f:cG�@�L�B�u�_�ø����#�f��ft �   #Ϻ������f��#�uf��ft@��f����t����뽋}3�������ك��E���8t3�����_�������������������������������������������������������������������������������������������U���0�E�E��M�Q�U��} t	�E�   ��E�    �E�E��}� u#h�uh�Yj j7h��j軳������u̃}� u0������    j j7h��h�h�u�Y������   �~  �} v	�E�   ��E�    �U�U�}� u#hvh�Yj j8h��j�@�������u̃}� u0�����    j j8h��h�hv��������   �  �   k� �E� �} ~�M�M���E�    �U��9Uv	�E�   ��E�    �E��E܃}� u#h �h�Yj j=h��j蜲������u̃}� u0������ "   j j=h��h�h ��:������"   �_  �} t	�E�   ��E�    �U؉Uԃ}� u#h��h�Yj j>h��j�!�������u̃}� u0�b����    j j>h��h�h���������   ��   �M��0�U����U��} ~A�E����t�U���EЋM����M���E�0   �U��EЈ�M����M��U���U빋E��  �} |>�M����5|3�E����E��M����9u�E�� 0�M����M���U�����M���U���1u�M�Q���E�P�&�M��Q�J�������P�U��R�EP蛹����3���]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���@���3ŉE��E�    �E�    �EP�M��˹���M�����Pj j j j �MQ�U�R�E�P�)����� �E�} t�M�UЉ�EP�M�Q�w������E�U��u8�}�u�E�   �M������E��j��}�u�E�   �M������E��N�:�E��t�E�   �M��u����E��0��M��t�E�   �M��W����E���E�    �M��C����E܋M�3��������]��������������������������������������������������������������������U��j �EP�MQ�������]����������U���@���3ŉE��E�    �E�    �EP�M��[����M�����Pj j j j �MQ�U�R�E�P������ �E�MQ�U�R�������E�E��u8�}�u�E�   �M��M����E��j��}�u�E�   �M��1����E��N�:�M��t�E�   �M������E��0��U��t�E�   �M�������E���E�    �M�������E��M�3�������]������������������������������������������������������������������U��j �EP�MQ�������]����������U��j �EP�MQ�UR������]����������������������U��j �EP�MQ�������]����������U���@���3ŉE��E�    �E�    �EP�M�諶���M������Pj j j j�MQ�U�R�E�P�	����� �E�MQ�U�R��������E�E��u8�}�u�E�   �M������E��j��}�u�E�   �M������E��N�:�M��t�E�   �M��c����E��0��U��t�E�   �M��E����E���E�    �M��1����E��M�3��������]������������������������������������������������������������������U��� �E�   �3�f�E��M�Q���  ��f�U��E�H�� �  f�M�U�B%�� �E�M��U��E��E�}� t�}��  t�P��  f�M��a�}� u)�}� u#�U�B    �E�     �Mf�U�f�Q�   �E�<  f�E��E�    ��M����  f�M��U����?  f�U��E���E�M�����U�B�E����M��U�B%   �uH�M���   �t	�E�   ��E�    �E�H��M��U�J�E���U�
f�E�f��f�E���M��U�ʋEf�H��]���������������������������������������������������������������������������������������������������U���,���3ŉE��EP�M�Q�:������U�Rj j���ċM���U�Pf�M�f�H�z������U�B�E֋M��UԋE�Pj jh��h �h8��M�Q�UR�EP������P�P������M�U�Q�E�M�3��2�����]������������������������������������������������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� ������������������������������������������������������SW3��D$�}G�T$���ڃ� �D$�T$�D$�}�T$���ڃ� �D$�T$�u�L$�D$3���D$���3�OyN�S�؋L$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$Oy���؃� _[� ���������������������������������������������̀�@s�� s����Ë�3������3�3������������������̀�@s�� s����Ë�3Ҁ����3�3�������������������U�� �]�������U���� ��E�M���u	�E�   ��E�    �U��U��}� u#h��h�Yj j*h�j谦������u̃}� u+������    j j*h�hx�h���N������E���M� ��E��]�������������������������������������������U����E%�����E�M#M��������   �} tj j �������U�3�t	�E�   ��E�    �M��M��}� u#h��h�Yj j,h��j�ȥ������u̃}� u-�	����    j j,h��hH�h���f������   �/�} t�EP�MQ�������U���EP�MQ�������3���]��������������������������������������������������������������U��j�˹����]������������������S�܃������U�k�l$���   ���3ŉE��C���h�����h�����t����C���x�����x�������x�����x���wR��x����$�d�ǅ|���   �Cǅ|���   �7ǅ|���   �+ǅ|���   �ǅ|���   ��K�   ǅ|���    ��|��� ��   ��t����P�K��Q��|���R��������u{�C��p�����p���t��p���t��p���t� �M����M��U������U��C�@�]��	�M�����M��S��R�C��P�KQ��|���R��t���P�M�Q�ܩ����h��  ��t����P�t�����ǅl���    �K�9t�=P� u�SR���������l�����l��� u�C�Q�������M�3��������]��[Ð��"�
����C�:�.���������������������������������������������������������������������������������������������������������������������������������������������U��3�]����������U��Q�E�    �E��U�+ȉM�u�M���t�E���E�M���M�σ}� }	�E�������}� ~�E�   �E���]����������������������������������U����E�E��M����tB�E�E��	�M����M��U����t�M���E��;�u
�E�+E����ыU����U�봋E�+E����]�����������������������������U��} u3��G�E���Et.�M���t$�E��U�;�u�M���M�U���U�ǋE� �M�+�]���������������������������U��Q�E���t=�U�U��	�E����E��M����t�E���U�;�u�E��֋M���M�3���]��������������������������������U���   ���3ŉE��E�H��  �U�JjU��P���P���������~Lj hj  h��h��h0���P���Q���������P��P���RjU�EP  P�ö����P�ڪ�����M�3��Ⱦ����]��������������������������������������������U����E�Q�s�������u	�E�   ��E�    �U�E��B�M�QR�F�������u	�E�   ��E�    �E�M��H�U�z t	�E�   ��E�Q�D  ���E�U�E�Bj jh��������M�Q��   t�E�H��   t�U�B��u
�M�A    ��]����������������������������������������������������������������U����E�Q�c�������u	�E�   ��E�    �U�E��B�M�y t	�E�   ��U�P�a   ���E��M�U��Qj jh����������E�H��u
�U�B    ��]�����������������������������������������U����E�    �} u3��X�Ef�f�M��U���U�E���A|	�M���Z~�U���a|'�E���z�M����M��Uf�f�E��M���M뾋E���]������������������������������U���   ���3ŉE������   ��x�����x����x tǅh���   �
ǅh���  j@��|���Q��h���R�EP�/�������u��x����A    �   ��  ��|���R��x����HQ�$��������  ��x����z tǅt���   �
ǅt���  j@��|���P��t���Q�UR赚������u��x����@    �   �S  ��|���Q��x����P諲������uf��x����Q��  ��x����Pj h�  h��h��h ��MQ���������P�URjU��x���P  P�ǲ����P�ަ�����&  ��x����Q���  ��x����x ��   ��x����QR��|���P��x����R�;�������ua��x����H����x����Jj h�  h��h��h ��EP�@�������P�MQjU��x�����P  R������P�2������}��x����H��uo�UR��  ����t_��x����H����x����Jj h�  h��h��h ��EP���������P�MQjU��x�����P  R蜱����P賥������x����H��   ��   �f  ��x����z tǅl���   �
ǅl���  h�   ��|���P��l���Q�UR薘������u��x����@    �   �4  ��|���Q��x����P茰��������  ��x����Q��   ��x����P��x����y ��   ��x����B   ��x����A�   k� ��x�����P  ��uJj h�  h��h��h ��EP��������P�MQjU��x�����P  R�b�����P�y������B  ��x����x ��   ��x����R�9�������x���;A��   ��x���Rj�EP�a  ����t|��x����Q��   ��x����P�   k� ��x�����P  ��uJj h�  h��h��h ��UR��������P�EPjU��x�����P  Q蘯����P诣�����{��x����B   ��x����A�   k� ��x�����P  ��uJj h�  h��h��h ��EP�@�������P�MQjU��x�����P  R������P�2�������x����H��uǅp���   �
ǅp���    ��p����M�3��������]� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE������   �����������x tǅ���   �
ǅ���  jx�����Q�����R�EP��������u������A    �   �   �����R������Q�u�������u_j hL  h��h��h ��UR�Ϳ������P�EPjU�������P  Q訬����P迠����������B��������A������B��uǅ ���   �
ǅ ���    �� ����M�3��n�����]� �������������������������������������������������������������������������������U��Q�} t�E���th���UR蠿������u5j�E�Ph  �M��P  Q��������u3��^�}� u��P�Kh���UR�V�������u'j�E�Ph   �M��P  Q�В������u3����UR裐�����E��E���]�������������������������������������������������U������3ŉE�j	�E�PjY�MQ�\�������u3��j	�UR�E�P��������u�   �3��M�3�������]������������������������U��V�EP��������u,�} t&�M�R����������E�Q������;�u3���   ^]�������������������������U����E�   �E�    �E�;Ed�}� t^�E�E�+����E�kM��U�
P�M�R萩�����E��}� ukE��M�T�E���}� }�M����M�	�U����U�딃}� u	�E�   ��E�    �E���]����������������������������������������������������U��������   �E��   k� 3ҋE�f��P  �M��A    �U�E���M���   �U��J�E��H���t�E���P�����Qh0��������U�����tw�U��B���t�U�R�j�������E�P�l������M��y uE�U�R�����Phh��i�������t'�M��Q���t�M�Q��������U�R��������E�P�@������M��y u3��  �} t�U��   �U���E�    �E�P�M�Q�E������E��}� t!�}���  t�}���  t�U�R� ��u3��G  �} t�E�M���} �*  �   k� 3ɋUf��   j h�   h��h �h8��E�P  P�ĺ������P�M���P  QjU�U��   R蜧����P賛����j@�EPh  �M��   Q�Վ������u3��   j@�U�   Rh  �E   P討������u3��vj_�M���   Q��������uj.�U�   R��������t'j@�E�   Pj�M��   Q�Q�������u3��j
j�U��   R�E�P��������   ��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���  ���3ŉE������   �������������  ������MQ�  ��������������z tǅ ���   �
ǅ ���  h�   �����P�� ���Q�����R�� ��u������     �   �   �����Q�������BP�ޤ������uD�����Q�  ����t1�����������B�����������Q��������������
��������uǅ����   �
ǅ����    �������M�3�������]� ������������������������������������������������������������������������������������U��������   �E��E��HQ�e�������u	�E�   ��E�    �U��E��Bjh0��� �M���u	�E�     ��]�����������������������������U��Q�E���  �U�
�� �E��E�M��H�U�E��B��]��������������U����Q����   �E��E��Q覶������u	�E�   ��E�    �U��E��B�M��QR�y�������u	�E�   ��E�    �E��M�H�U�B    �E��x t	�E�   ��M��R�M  ���E��E��M��Hjh��� �U�%   t�M���   t
�E���u	�U�    ��]������������������������������������������������������������������U����1����   �E��E��Q膵������u	�E�   ��E�    �U��E��B�M��y t	�E�   ��U��P�d   ���E�M��U�Qjh���� �E���u	�U�    ��]��������������������������������������������������U����E�    �Ef�f�M��U���U�E���A|	�M���Z~�U���a|'�E���z�M����M��Uf�f�E��M���M뾋E���]����������������������������������������U���  ���3ŉE��Լ���   ������ļ�����  ������MQ��  ���� ���������z tǅ����   �
ǅ����  h�   �����P������Q�� ���R�� ��u������     �   ��  �����Q������BP����������  ������y tǅ����   �
ǅ����  h�   �����R������P�� ���Q�� ��u������    �   �k  �����P������R袟������u9��������  ������
������� ����H������� ����B��   ����������   ������x tu������QR�����P������R�d�������uO��������������
������� ����H������P�m����������;Au������� ����B�B��������u5�� ���P�q  ����t"��������������������� ����Q��������   ��   ��  ������z tǅ����   �
ǅ����  h�   �����P������Q�� ���R�� ��u������     �   ��  �����Q������P���������  ��������   ������������y t5������   ������������z u������� ����H�   ������z tj������Q�����������;BuN�����Pj�� ���Q�~  ����t0������   ������������z u������� ����H�0������   ������������z u������� ����H�   ������z uu������x ti�����Q������P�ɜ������uM�����Qj �� ���R��  ����t1��������   ������
������x u������� ����Q��������uǅ����   �
ǅ����    �������M�3��դ����]� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���  ���3ŉE������   �� ����������  ������MQ�  ��������� ����z tǅ����   �
ǅ����  h�   �����P������Q�����R�� ��u������     �   �$  �����Q�� ����P�_�������u^�� ����y u�����Rj�����P�Q  ����t1�����������Q�����������H���������������   �� ����z uu�� ����x ti�����Q�� ����P�͙������uM�����Qj �����R��  ����t1�����������H�����������B����������������������uǅ����   �
ǅ����    �������M�3��١����]� ��������������������������������������������������������������������������������������������������������������������������U����E�    �Ef�f�M��U��U�E���E�}� tO�M���a|�U���f�E���'f�E���M���A|�U���F�E���f�E��M����U��DЉE�둋E���]����������������������������������������������U��Q�} t�E���th���UR�0�������u0j�E�Ph  �M�QR�� ��u3��Y�}� u��K�Fh���EP��������u"j�M�Qh   �U�BP�� ��u3����MQ�=}�����E��E���]�������������������������������������������U���f�Ef�E��E�    �	�M����M��}�
s�U��E��E��;�u3���ظ   ��]�������������������������U���V�E%�  �ȁ�   �щU��ز���   �E�j�E�Ph   �M�Q�� ��u3��9�U;U�t,�} t&�E��Q���������U��P������;�u3���   ^��]������������������������������������������U����E�   �E�    �E�;Ed�}� t^�E�E�+����E�kM��U�
P�M�R�������E��}� ukE��M�T�E���}� }�M����M�	�U����U�딃}� u	�E�   ��E�    �E���]����������������������������������������������������U���$���3ŉE��g����   �E�jj �E�P�������J����  �E܋M܍U���E܋�M�} u�U�R�������(  �E�M��U�   �E�P�M�y t*�U�B���t�U��R�����Ph0��������M��    �U�: ��   �E������   �E�x t�M�Q���t�M�Q�1�������U�R�C������E�8 uO�M�Q�����Rhh���������t0�E�x t�M�Q���t�M�Q���������U�R��������0�E�x t�M�Q���t�M�Q���������U�R�Z������E�8 u3��!  �} t�M��   �M���E�    �U�R�E�P�������E�}� t!�}���  t�}���  t�M�Q� ��u3���   j�U�BP�� ��u3��   �} t�M�U�jU�E�P  P�M�QR董�����} txjU�E   P�M�QR�q�����j@�EPh  �M�QR�� ��u3��Cj@�E�   Ph  �M�QR�� ��u3��j
j�E   P�M�Q�U������   �M�3��6�����]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E������E�    �E�    �} t	�E�   ��E�    �E؉Eԃ}� u#h��h�Yj jmh�j�${������u̃}� u.�e����    j jmh�ht�h���¹���������   �U�U��E����E��M��Q��U��E�    �E�    j �E�Pj@�MQ�UR�E�P�M�Q�ϋ�����E��E������   �Q�}� tJ�}� t8�U����E������0��T����E����M������0��T�M�Q�x����Ã}� t�����U܉�����E�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������U����E�    �E������E�E��M����M��U��B��E��E�    j �M�Q�U�R�EP�MQ�UR�������E�}� t	�E�������E�E��E���]���������������������������������U��j�hx�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�   ��E�    �E��E܃}� u&h��h�Yj h�   h�j�x������u̃}� u3�����    j h�   h�h��h���:������   ��  �U������} t	�E�   ��E�    �E؉Eԃ}� u&h��h�Yj h�   h�j�x������u̃}� u3�V����    j h�   h�h��h��谶�����   �9  �} ��   �U�����u	�E�   ��E�    �EЉẼ}� u&h��h�Yj h�   h�j�w������u̃}� u3�ƽ���    j h�   h�h��h��� ������   �   �E�    �UR�EP�MQ�UR�EP�MQ�U�R�F������E��E������   �[�}� tT�}� t@�E����U�������0��T����E����E� ������0��T�U�P�{t����Ã}� t	�M������E�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    �E�P�MQ��������u����8�U R�EP�MQ�UR�E�P�MQ�UR�@z�����E�j�E�P�%������E���]�������������������������������U��j�EP�MQ�UR�EP�MQ������]��������������U��j �EP�MQ�UR�ƃ����]����������������������U���T�} u3���  �EP�M��~���M�������H�y u'�UR�EP�MQ�
������EԍM�������E��  �} t	�E�   ��E�    �U�U��}� u#h8�h�Yj j>hX�j�it������u̃}� u=誺���    j j>hX�h��h8��������E�����M��8����E��2  �} t	�E�   ��E�    �M�M�}� u#h��h�Yj j?hX�j��s������u̃}� u=�"����    j j?hX�h��h���������E�����M�谍���E��  �E�EȋM���M�}� �  �Uf�f�E��M���M�M��w����P�E��L��t|�} u@3�f�U��M��R����@�M��D��t	�E�    �	�M��U�f�E�f�E��   �M���u	�E�    ��E����M�E��E���Ef�M�f�M��Uf�f�E��M���M�M��ο���P�E��L��tM�} u3�f�U��?�E���E�M���u	�E�    ��E����M�E܋E���Ef�M�f�M��U��E�;�t/�M��U�;�~	�E�   ��E������E؉EčM��6����E��3�M���u�E�    �M������E���h����E�    �M������E���]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR������]����������������������U���XV�EP�M��z���} u�E�    �M��׊���E��	  �M��˽���H�y u'�UR�EP�MQ�������EЍM�蟊���E���  �} t	�E�   ��E�    �U�U��}� u#h8�h�Yj j?h �j�Hp������u̃}� u=艶���    j j?h �hl�h8��������E�����M������E��I  �} t	�E�   ��E�    �M�M�}� u#h��h�Yj j@h �j��o������u̃}� u=�����    j j@h �hl�h���^������E�����M�菉���E���  �E�EċM���M�}� ��  �Uf�f�E��M���M�M��V����P�E��L���>  �} u@3�f�U��M��-����@�M��D��t	�E�    �	�M��U�f�E�f�E���  �M���u3�f�E���   �M����U��f�M��M���M�u��M�辻���P�   k� �T
;�|C�u��M�螻���@�   �� �T;�#�M�肻���@�   ���T�E��f�E��b�u��M��[����H�   k��L;�|B�u��M��;����P�   ���L;�"�M������P�   k��T
�E��f�E��D�M�������H�U��D��t�M������H�U���  �E���M��M�f�U�f�U��Ef�f�M��U���U�M�裺���@�M��T���  �} u3�f�E��E  �M���M�U���u3�f�M���   �U����E��f�U��U���U�u��M��7����@�   k� �D;�|C�u��M������H�   �� �D;�#�M�������H�   ���D�M��f�M��b�u��M��Թ���P�   k��T
;�|B�u��M�费���@�   ���T;�"�M�蘹���@�   k��D�M��f�M��D�M��t����P�E��L��t�M��[����P�E���  �M���U��U�f�E�f�E��M��U�;�t/�E��M�;�~	�E�   ��E������U؉U��M�������E��3�E���u�E�    �M������E���Q����E�    �M��Ʌ���E�^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U�����n����teh��h@��� P�� �E��}� u����c�E�   �E�E�M �M��E�    �U�U��E�    �E�P�MQ�UR�EP�MQ�U��#j �UU R�EP�MQ�UR�EP�MQ�T��]������������������������������������������������������U��j�h،h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E������E�    �E�    �} t	�E�   ��E�    �E؉Eԃ}� u#h��h�Yj jmh�j�i������u̃}� u.�E����    j jmh�h��h��袧���������   �U�U��E����E��M��Q��U��E�    �E�    j �E�Pj@�MQ�UR�E�P�M�Q�/m�����E��E������   �Q�}� tJ�}� t8�U����E������0��T����E����M������0��T�M�Q��e����Ã}� t�i����U܉�����E�M�d�    Y_^[��]����������������������������������������������������������������������������������������������������������U����E�    �E������E�E��M����M��U��B��E��E�    j �M�Q�U�R�EP�MQ�UR�������E�}� t	�E�������E�E��E���]���������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �E�    �} t	�E�   ��E�    �E��E܃}� u&h��h�Yj h�   h�j�f������u̃}� u3������    j h�   h�h��h���������   ��  �U������} t	�E�   ��E�    �E؉Eԃ}� u&h��h�Yj h�   h�j��e������u̃}� u3�6����    j h�   h�h��h��萤�����   �9  �} ��   �U�����u	�E�   ��E�    �EЉẼ}� u&h��h�Yj h�   h�j�ee������u̃}� u3覫���    j h�   h�h��h��� ������   �   �E�    �UR�EP�MQ�UR�EP�MQ�U�R�i�����E��E������   �[�}� tT�}� t@�E����U�������0��T����E����E� ������0��T�U�P�[b����Ã}� t	�M������E�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   �E�    �E�    �E�    �E� �E�    ǅ`���   ǅd���    �E%�   tǅh���    �E��ǅh���   �E� j h:  h�h��h���M�Q�g�����P�n�����U�� �  u/�E% @ t�M��ɀ   �M���}� �  t�U��ʀ   �U��E���E�t�}�t�}�t6�@�E�   ���   �M��t�U��   t	�E�   ���E�   @�   �E�   ��   ��g���     �E� ����3�t	�E�   ��E�    �U��U��}� u&h$�h�Yj ha  h�j�Hb������u̃}� u3艨���    j ha  h�h��h$��������   �  �M�M��U����U��}�pw_�E������$����E�    ��   �E�   ��   �E�   ��   �E�   �   �}�   �u	�E�   ��E�    �   ��f���     �U�����3�t	�E�   ��E�    �M���x�����x��� u&hh�h�Yj h�  h�j�;a������u̃�x��� u3�y����    j h�  h�h��hh��ӟ�����   �   �E%   �E�}�   7�}�   tK�}�   �}�   t]�}� t3�}�   t6�d�}�   tO�Y�}�   t,�}�   t/�}�   t�<�E�   ��   �E�   ��   �E�   �   �E�   �   �E�   �   �e���     �M�����3�tǅ|���   �
ǅ|���    ��|�����l�����l��� u&h$�h�Yj h�  h�j��_������u̃�l��� u3�0����    j h�  h�h��h$�芞�����   �  �EȀ   �E�    �U��   t�����#E%�   u�E�   �M��@t �U���   �U��E�   �E��M����M��U��   t�E�   �EȋM��    t�U���   �U��E�� t�M���   �M���U��t�E�   �E���z���M��U�:�u+�7d���     �E� �����(����    ����� ��
  �M�   �U�R�E�P�M�Q��`���R�E�P�M�Q�UR�8������E�}���  �E�%   �=   ���   �M����   �U�������U��E�P�M�Q�U�R��`���P�M�Q�U�R�EP��������E�}��u^�M����E�������0��D
����M����M�	������0��D
�� P�\�����*���� �E���	  �^�M����E�������0��D
����M����M�	������0��D
�� P�Q\�����ʣ��� �E��r	  �M�Q�� �E��}� ��   �E�    �U����M�������0��L����U����U�������0��L�� �E��M�Q��[�����U�R�� �}� u�8����    �-���� �E���  �}�u�M���@�M���}�u
�U����U��E�P�M�R�#|�����E����E��M����E�������0��E��D
�M����E�������0��D
$$��M����M�	������0��D
$�E���H�  �M���   �  �U����   jj�j��E�Q�4������EЉUԋU�#Uԃ��u/�.a���8�   t�E�Q賌����������U���  �   3�f�E�j�M�Q�U�P�{������uA�M���u8�U�R�E�P�M�R�!��������u�E�Q�O�����贡����U��\  j j j �E�Q聂�����EЉUԋU�#Uԃ��u�E�Q�������r�����U��  �E�%�   �  �M�� @ u'�U��� @ u�E @  �E��M��� @ M�M�U�� @ u&h��h�Yj h�  h�j�Z������u̋M�� @ �M؁}�   &�}�   tW�}� @  t1�}�   t.�}� @ t%�D�}� @ t1�}�   t.�}� @ t%�'�E� �!�U��  ��  u�E��
�E���E��E%   �&  �E�    �E�    �E�    �M���@��  �U���   ��U��}�   @t'�}�   �t�}�   ���   �q  �E�   �e  �E�E��M����M��}���   �U��$�(�jj j �E�Q迀������X�����\�����X����\���tPj j j �E�Q葀������@�����D�����@���#�D������u�E�Q�������v�����U��  ��E�   �   �E�E��M����M��}���   �U��$�<�jj j �E�Q��������H�����L�����H����L���tWj j j �E�Q��������P�����T�����P���#�T������u�E�Q�d������ɞ����U��q  �E�   ��E�   ��E�   �}� ��  j�E�P�M�R�Cx������p�����p��� ~7�}�u13�u&hL�h�Yj h�  h�j��W������u��E�    ��p����U��}��t�}�t:�}�t"��   �E�Q誈����������U��  �}�﻿ u	�E���   �E�%��  =��  uO�M�R�l�����3�u&h��h�Yj h  h�j�`W������u�觝���    �E�   �G  �U܁���  ����  uHj j j�E�Q�[~�����EЉUԋU�#Uԃ��u�E�Q�������L�����U���  �E��Bj j j �E�Q�~�����EЉUԋU�#Uԃ��u�E�Q蟇����������U��  �}� ��   �E�    �E�    �E�    �E���t�����t���t��t���t��E���  �E�   ��E�﻿ �E�   �M�;M�~U�E�    �U�+U�R�EčL�Q�U�P�{�����E��}��u�M�R�������X���� �E��   �M�M��M�룋U����M�������0��M����T$��
ыE����E� ������0��T$�U��   u	�E�    ��E�   �E����U�������0��U������D$$
M����M�	������0��D
$�E���HuH�M��t@�U����M�������0��L�� �U����U�������0��L�M���   ���   ���   �U����   �E�P�� �M�������M��E�   �U�R�E�P�M�Q��`���R�E�P�M�Q�UR�4������E�}��uk�� P�LS�����E����U�������0��T����E����E� ������0��T�U�P�p�����w�����M��"� �U����M�������0��M��E��]Ë������������� �I w�w�����w�4�4�����4�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�EP�MQ�UR�EP�MQ�݃����]��������������U���$�=� ��  �E�    �} ��  �} t	�E�   ��E�    �E�E��}� u#h�h�Yj jmh@�j�N������u̃}� u0�͔���    j jmh@�h��h��*����������D  �} t	�E�   ��E�    �U�U�}� u#h��h�Yj jnh@�j�N������u̃}� u0�R����    j jnh@�h��h��诌����������   �M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���M�U���U�E���Et�M���t�U��E�;��a����M��U�+ʉM܋E���j �EP�MQ�UR�}������]��������������������������������������������������������������������������������������������������������������������������U���4�E�    �} �@  �} t	�E�   ��E�    �E�E��}� u#h�h�Yj j=h@�j�9L������u̃}� u0�z����    j j=h@�h��h��׊����������  �} t	�E�   ��E�    �U�U�}� u#h��h�Yj j>h@�j�K������u̃}� u0������    j j>h@�h��h���\����������M  �MQ�M��<U���M�肘����   �����    ��   �M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���A|�E���Z�U��� �E��	�M��U�f�E�f�E��M���M�U���U�E���Et�M���t�U��E�;��a����i�M����P�M�R��G����f�E��M�覗��P�E�Q��G����f�E��U���U�E���E�M���Mt�U���t�E��M�;�t��U��E�+ЉU܍M��Hd���E܋�]�������������������������������������������������������������������������������������������������������������������������������������������������������������������U���x  ���3ŉE�ǅ(���    ǅ����    ǅx���    ǅ����    ǅT���    ǅ���    ǅ4���    ǅ����    ǅ@���    �EP��`�����R��ǅ����    ǅp���    ǅ����    ǅ����    ǅ��������ǅ��������ǅ|�������ǅ��������ǅ��������ǅH���    ������������} tǅ����   �
ǅ����    ������������������ u&h �h�Yj h  hx�j�SH������u̃����� uI葎���    j h  hx�h��h �������ǅx���������`����b����x����1;  �E�������������Q��@��   ������P�H{������\�����\����t-��\����t$��\�������\��������0��������
ǅ������������H$�����х�uV��\����t-��\����t$��\�������\��������0��������
ǅ������������B$�� ���ȅ�tǅ����    �
ǅ����   ������������������ u&hp�h�Yj h	  hx�j��F������u̃����� uI�����    j h	  hx�h��hp��n�����ǅ����������`����`���������9  �} tǅ����   �
ǅ����    ������������������ u&h��h�Yj h  hx�j�-F������u̃����� uI�k����    j h  hx�h��h���ń����ǅ����������`�����_���������9  ǅ����    �E������ǅ����    �����������������������8  ������u������ u�8  ǅ����    ǅX���    ǅH���    ǅ ���    ǅ��������ǅx���    ǅ����    �������Uǅ��������ǅ|�������ǅ��������ǅ���������E��������������������E���E������ �5  ������ ��4  �������� |%��������x��������(����������
ǅ����    ������������k�����	��X�����H�����X�����X�����  �E���%��  �������u\j
��p���R�EP�n������~9��p������$u+������ uh@  j ������P�k����ǅ����   �
ǅ����    �������.  j
��p���Q�UR�Nn��������������p������E������ ��   ������ |#��p������$u������d}ǅ����   �
ǅ����    ������������������ u&h�h�Yj hU  hx�j�<C������u̃����� uI�z����    j hU  hx�h��h��ԁ����ǅ����������`�����\���������6  ������;�����~��������������������������������������   ��X�����   3�tǅ����   �
ǅ����    ������������������ u&h��h�Yj ha  hx�j�OB������u̃����� uI荈���    j ha  hx�h��h��������ǅ����������`����\���������-5  ��X����������������2  �������$�������� u	������t������u�������u��1  ǅ@���    ��`���觎��P������R趏��������   ������P�MQ������R�#I  ���E��������U���U��������tǅ����   �
ǅ����    ������������������ u&h�h�Yj h�  hx�j��@������u̃����� uI�3����    j h�  hx�h��h������ǅ����������`����Z����������3  ������P�MQ������R�FH  ���0  ǅ���    �������4�����4�����x�����x�����T���ǅ����    ǅ��������ǅ@���    �O0  ��������$�����$����� ��$�����$���wj��$������$�����������������E���������������4���������������#�������ɀ   ����������������������/  ��������*��  ������ u�MQ�MV������x����  j
��p���R�EP��i��������|�����p������M������ �'  ��|��� |#��p������$u������d}ǅ����   �
ǅ����    ������������������ u&h �h�Yj h�  hx�j��>������u̃����� uI�����    j h�  hx�h��h ��^}����ǅp���������`����X����p����1  ��|���;�����~��|������������������������������������|����������� uE��|�����Ǆ����   ��|�������������������|�������������������   ������Q������Rj��|�����������Q�o������tǅ����   �
ǅ����    ������������������ u&h��h�Yj h�  hx�j�i=������u̃����� uI觃���    j h�  hx�h��h���|����ǅ����������`����,W���������G0  �/-  �+��|�������������h�����h���P�S������x�����x��� }����������������x����ډ�x����k�x���
�������TЉ�x����,  ǅ����    �,  ��������*��  ������ u�MQ�@S�����������  j
��p���R�EP��f��������������p������M������ �'  ������ |#��p������$u������d}ǅ���   �
ǅ���    ����������������� u&h��h�Yj h�  hx�j�;������u̃����� uI������    j h�  hx�h��h���Qz����ǅ����������`����|U���������.  ������;�����~��������������������������������������������������� uE��������Ǆ����   ������������������������������������������   ������Q������Rj��������������Q�l������tǅ����   �
ǅ����    ���������������� u&h8�h�Yj h�  hx�j�\:������u̃���� uI蚀���    j h�  hx�h��h8���x����ǅ`���������`����T����`����:-  �"*  �+��������������������������P�P���������������� }
ǅ���������k�����
�������DЉ�������)  ������������������I����������.�B  �������4�$� �U���lu�M���M��������   �����������������������   �M���6u+�E�H��4u�U���U������ �  �������   �M���3u(�E�H��2u�U���U������%����������e�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu��������   �������ǅX���    �����"�������� �������������   �������S(  �������� ����� �����A�� ����� ���7��%  �� �������$�d��������0  u������   ��������������  ��  ǅt���    ������ u�UR��s����f��,����  ������ |������d}ǅ����   �
ǅ����    ������������������ u&h��h�Yj h�  hx�j�:7������u̃����� uI�x}���    j h�  hx�h��h����u����ǅX���������`�����P����X����*  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R�?h������tǅ|���   �
ǅ|���    ��|��������������� u&h@�h�Yj h�  hx�j�6������u̃����� uI�B|���    j h�  hx�h��h@��t����ǅ����������`�����O����������(  � #  �,����������������P�����P���Q��q����f��,�����,���Rh   ������P������Q��|������t�����t��� t
ǅ4���   �^  ������ u�UR��K����f��8����  ������ |������d}ǅ����   �
ǅ����    ��������l�����l��� u&h��h�Yj h�  hx�j�4������u̃�l��� uI��z���    j h�  hx�h��h���Rs����ǅ����������`����}N���������'  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R�e������tǅ����   �
ǅ����    ��������d�����d��� u&h��h�Yj h�  hx�j�3������u̃�d��� uI��y���    j h�  hx�h��h���r����ǅH���������`����GM����H����b&  �   �,��������������������������Q��I����f��8����   k� ��8���������ǅ����   �������������B   ������ u�EP�I������D����  ������ |������d}ǅ����   �
ǅ����    ��������\�����\��� u&h��h�Yj h�  hx�j�L2������u̃�\��� uI�x���    j h�  hx�h��h����p����ǅ@���������`����L����@����*%  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������P������Qj��������������P�Qc������tǅ����   �
ǅ����    ��������T�����T��� u&h��h�Yj h�  hx�j�1������u̃�T��� uI�Tw���    j h�  hx�h��h���o����ǅ����������`�����J����������#  �2  �+����������������8�����8���R�lG������D�����D��� t��D����x u#�p�������������R�Z�����������d������%   t/��D����Q��������D���� �+���������ǅ@���   �(ǅ@���    ��D����Q��������D�����������d  ��������0  u������   �������������uǅ����������������������������<��������� u�EP�dF�����������  ������ |������d}ǅL���   �
ǅL���    ��L��������������� u&h��h�Yj h:  hx�j�"/������u̃����� uI�`u���    j h:  hx�h��h���m����ǅ����������`�����H��������� "  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������P������Qj��������������P�'`������tǅD���   �
ǅD���    ��D��������������� u&h��h�Yj h>  hx�j��-������u̃����� uI�*t���    j h>  hx�h��h���l����ǅ0���������`����G����0�����   �  �+��������������������������R�BD����������������%  ��   ������ u�t�������ǅ@���   �������������<�����(�����<�������<�����(��� t��������t������������뾋����+��������������t������ u�p��������������������<�����������<�������<��������� t��������t������������뾋����+�������������  ������ u�UR�C�����������  ������ |������d}ǅ<���   �
ǅ<���    ��<��������������� u&h��h�Yj h�  hx�j��+������u̃����� uI�r���    j h�  hx�h��h���pj����ǅ ���������`����E���� ����  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R��\������tǅ4���   �
ǅ4���    ��4��������������� u&h��h�Yj h�  hx�j�*������u̃����� uI��p���    j h�  hx�h��h���:i����ǅ����������`����eD���������  �  �+������������������������Q��@������������a������   3�tǅ,���   �
ǅ,���    ��,��������������� u&h�h�Yj h�  hx�j�)������u̃����� uI��o���    j h�  hx�h��h��Th����ǅ����������`����C���������  ��  �������� t������f������f���������������ǅ4���   �  ǅ���   �������� ��������������@��������������  ������ ��  ������ |������d}ǅ$���   �
ǅ$���    ��$��������������� u&h��h�Yj h�  hx�j�(������u̃����� uI��n���    j h�  hx�h��h���g����ǅ���������`����HB��������c  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R�Y������tǅ���   �
ǅ���    ����������������� u&h(�h�Yj h�  hx�j�\'������u̃����� uI�m���    j h�  hx�h��h(���e����ǅ����������`����A���������:  �x  ������������ǅ ���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Yh�  hp�j��������]  Q�"������H�����H��� t��H���������������]  �� ����
ǅ�����   ������ u#�M���M�U�B��J���|����������!  ������ |������d}ǅ���   �
ǅ���    ����������������� u&h��h�Yj h  hx�j�%������u̃����� uI��k���    j h  hx�h��h���Gd����ǅ���������`����r?��������  ������t&h��h�Yj h  hx�j�.%������u̋������������������������������������B��J���|�����������`�����q��P�����R������P������Q�� ���R������P��|���Q�   k���0�Q� �Ѓ���������   t6������ u-��`����q��P������P�   k�	��0�P� �Ѓ���������gu;��������   u-��`����Eq��P������P�   ����0�R� �Ѓ����������-u!��������   ��������������������������Q�N�����������?  ��������@������ǅ0���
   �   ǅ0���
   �   ǅ����   ǅ(���   �
ǅ(���'   ǅ0���   ������%�   t2�   k� Ƅt���0��(�����Q�   �� ��t���ǅT���   �)ǅ0���   ��������   t������   �������������� �  �N  ������ u�UR�R�����������������#  ������ |������d}ǅ����   �
ǅ����    ������������������ u&h��h�Yj h�  hx�j�p"������u̃����� uI�h���    j h�  hx�h��h���a����ǅ����������`����3<���������N  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R�uS������tǅ����   �
ǅ����    ������������������ u&h�h�Yj h�  hx�j�:!������u̃����� uI�xg���    j h�  hx�h��h���_����ǅ ���������`�����:���� ����  �V  �1����������������t�����t���Q��O������������������  ��������   �N  ������ u�EP�O�����������������#  ������ |������d}ǅ����   �
ǅ����    ��������x�����x��� u&h��h�Yj h�  hx�j� ������u̃�x��� uI�Nf���    j h�  hx�h��h���^����ǅl���������`�����9����l�����  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������P������Qj��������������P�Q������tǅp���   �
ǅp���    ��p�����h�����h��� u&h��h�Yj h�  hx�j��������u̃�h��� uI�e���    j h�  hx�h��h���r]����ǅd���������`����8����d����  ��  �1����������������\�����\���R�|M�����������������r	  �������� ��  ��������@�R  ������ u�UR��4�������������������%  ������ |������d}ǅ`���   �
ǅ`���    ��`�����X�����X��� u&h��h�Yj h�  hx�j�������u̃�X��� uI��c���    j h�  hx�h��h���:\����ǅT���������`����e7����T����  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R�N������tǅP���   �
ǅP���    ��P�����H�����H��� u&h��h�Yj h�  hx�j�l������u̃�H��� uI�b���    j h�  hx�h��h���[����ǅL���������`����/6����L����J  �	  �3����������������D�����D���Q��2�������������������Q  ������ u!�UR�2��������������������'  ������ |������d}ǅ@���   �
ǅ@���    ��@�����8�����8��� u&h��h�Yj h�  hx�j�N������u̃�8��� uI�a���    j h�  hx�h��h����Y����ǅ<���������`����5����<����,  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������R������Pj��������������R�SL������tǅ0���   �
ǅ0���    ��0�����(�����(��� u&h��h�Yj h  hx�j�������u̃�(��� uI�V`���    j h  hx�h��h���X����ǅ4���������`�����3����4�����  �4  �5����������������,�����,���Q�n0��������������������  ��������@�P  ������ u�EP�50������������������$  ������ |������d}ǅ ���   �
ǅ ���    �� ������������� u&h��h�Yj h  hx�j��������u̃���� uI�*_���    j h  hx�h��h���W����ǅ$���������`����2����$�����  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������P������Qj��������������P��I������tǅ���   �
ǅ���    ��������������� u&h��h�Yj h  hx�j�������u̃���� uI��]���    j h  hx�h��h���NV����ǅ���������`����y1��������
  ��  �2������������������������R�.������������������M  ������ u�EP��-����3ɉ������������%  ������ |������d}ǅ ���   �
ǅ ���    �� ��������������� u&h��h�Yj h4  hx�j�������u̃����� uI��\���    j h4  hx�h��h���3U����ǅ���������`����^0��������y	  ������ �0  �������������� uE��������Ǆ����   ������������������������������������������   ������Q������Rj��������������Q�G������tǅ����   �
ǅ����    ������������������ u&h��h�Yj h8  hx�j�e������u̃����� uI�[���    j h8  hx�h��h����S����ǅ���������`����(/��������C  �  �3��������������������������P�+����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�L�����P�����������   ���������������L�����������P����������� �  u(������%   u��L�����P����� ��L�����P��������� }ǅ����   �%���������������������   ~
ǅ����   ��L����P���u
ǅT���    �   i��  �������������������������������������������� ��L����P�����   ��0����RP��P���R��L���P�
-����0�������0����RP��P���Q��L���R�F+����L�����P��������9~������(�����������������������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0��������������������u������ u�  ��4��� �b  ��������@tv��������   t�   k� Ƅt���-ǅT���   �L��������t�   k� Ƅt���+ǅT���   �%��������t�   k� Ƅt��� ǅT���   ��x���+�����+�T�����������������u������Q�UR������Pj �7  ��������Q������R�EP��T���Q��t���R�_  ����������t'��������u������R�EP������Qj0��  ����@��� ��   ������ ��   ǅ����    �������������������������������������������������������� ��   ������f�f������������Rj�E�P������Q�>X������������������������������ u	������ uǅ���������*������P������Q�UR������P�M�Q�D  ���N����(������R������P�MQ������R������P�  �������� |'��������t������R�EP������Qj �  ����H��� tj��H���R�����ǅH���    �������X��� t��X���tǅ����    �
ǅ����   ������������������ u&hh�h�Yj h�  hx�j�{������u̃����� uI�U���    j h�  hx�h��hh��N����ǅ����������`����>)���������Y  �������*  ������ �  ǅ����    ���������������������;�������  �������������������������������������  ������$�����������E�������MQ�X%�����  ���������E�������MQ�J�����d  ���������E�������MQ�%�����@  ���������E�������MQ�8=�����  ���������E�������MQ�=������   ���������E�������MQ�$������   ���������E�������MQ�\�����������������   3�tǅ����   �
ǅ����    ������������������ u&h��h�Yj h2	  hx�j�F������u̃����� uF�S���    j h2	  hx�h��h����K����ǅ����������`����	'���������'������1�����������������`�����&���������M�3��+����]Ð���c��������_������������� �I h�8�,�I�Z� �j����� �������:�a����   	
�:^��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���<�E�    �E�    �E�H��pt	�U��pu'�E�H�U;�u	�E�   ��E�    �E��  �E�H��st�U�B��St	�E�    ��E�   �M��M��U��st�E��St	�E�    ��E�   �M�M��}� u�}� ta�U�;U�uJ�E�H��  t	�E�   ��E�    �U��  t	�E�   ��E�    �E�;E�u	�E�   ��E�    �E���  �M�Q��dtv�E�H��itj�U�B��ot^�M�Q��utR�E�H��xtF�U�B��Xt:�M��dt1�U��it(�E��ot�M��ut�U��xt�E��X�,  �M�Q��dtE�E�H��it9�U�B��ot-�M�Q��ut!�E�H��xt�U�B��Xt	�E�    ��E�   �M��dt6�U��it-�E��ot$�M��ut�U��xt�E��Xt	�E�    ��E�   �M�;M�t3��   �U�B%   t	�E�   ��E�    �M��   t	�E�   ��E�    �U�;U�u;�E�H�� t	�E�   ��E�    �U�� t	�E�   ��E�    �E�;E�t3���M�;Uu	�E�   ��E�    �Eċ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E����U�
�E��A��Q�]��������������������U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�7�����E��}��u�M�������U����M���]�������������������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��|�U�    �E�E��M���M�}� ~N�U��E��MQ�UR�E�P�w������M���M�U�:�u�E�8*u�MQ�URj?�L�������띋E�8 u�M�U���]������������������������������������������������U���P  ���3ŉE�ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    �EP��P�������ǅ����    �<����p����} tǅD���   �
ǅD���    ��D������������� u&h �h�Yj h  hx�j�]�������u̃���� uI�;���    j h  hx�h��h ���3����ǅ����������P���� ���������  �E�� ����� ����Q��@��   �� ���P�R(�����������������t-�������t$�������������������0��������
ǅ������������H$�����х�uV�������t-�������t$�������������������0��������
ǅ������������B$�� ���ȅ�tǅL���    �
ǅL���   ��L������������� u&hp�h�Yj h	  hx�j���������u̃���� uI�:���    j h	  hx�h��hp��x2����ǅ����������P�������������A  �} tǅ���   �
ǅ���    �������<�����<��� u&h��h�Yj h  hx�j�7�������u̃�<��� uI�u9���    j h  hx�h��h����1����ǅ����������P��������������  ǅ����    ǅ����    ǅ����    ǅ����    ǅ|���    �E��������������������E���E������ �i  ������ �\  �������� |%��������x��������(���������
ǅ���    �����������k�����	��������H�����������������   3�tǅ4���   �
ǅ4���    ��4��������������� u&h��h�Yj he  hx�j��������u̃����� uI��7���    j he  hx�h��h���I0����ǅ����������P����t���������  ��������,�����,����%  ��,����$�XFǅ����    ��P����2>��P������R�A?��������   ������P�MQ������R�  ���E��������U���U��������tǅ���   �
ǅ���    �������$�����$��� u&h�h�Yj h�  hx�j��������u̃�$��� uI�6���    j h�  hx�h��h��/����ǅ����������P����C
����������  ������P�MQ������R��  ����  ǅ����    ������������������������������������ǅ����    ǅ��������ǅ����    �  �������������������� ������������wj���������F�$�xF���������������E���������������4���������������#�������ɀ   ����������������������  ��������*u:�MQ������������������ }���������������������؉������k�����
�������DЉ������  ǅ����    �  ��������*u'�UR�s���������������� }
ǅ���������k�����
�������TЉ������F  ��������������������I������������.�3  ���������F�$��F�M���lu�E���E��������   �����������������������   �E���6u,�U�B��4u �M���M�������� �  �������   �E���3u)�U�B��2u�M���M������������������S�E���dt7�U���it,�M���ot!�E���ut�U���xt�M���Xu�ǅ����    ������#�������� ���������������   ��������  ��������������������A������������7�)
  ��������$G�$��F������%0  u��������   ��������������  t[ǅ����    �EP��(����f��t�����t���Qh   ������R������P��3���������������� t
ǅ����   �2�MQ�	����f��l����   k� ��l���������ǅ����   �������������J	  �EP������������������ t�������y u#�p�������������P�������������e��������   t/�������B��������������+���������ǅ����   �(ǅ����    �������B��������������������  ������%0  u��������   �������������uǅ������������������������������MQ��������������������  ��   ������ u�t�������ǅ����   �������������������������������������������� t���������t��������������뾋�����+��������������u������ u�p��������������������������������������������������� t���������t��������������뾋�����+������������*  �MQ� ������8����!������   3�tǅH���   �
ǅH���    ��H�����@�����@��� u&h�h�Yj h�  hx�j�j�������u̃�@��� uI�/���    j h�  hx�h��h��(����ǅ����������P����-����������	  �_  �������� t��8���f������f����8����������ǅ����   �%  ǅ����   �������� ��������������@������������������ǅ|���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Zh�  hp�j��������]  R�=����������������� t ��������������������]  ��|����
ǅ�����   �U���U�E�H��P���������������P�����4��P������P������Q������R��|���P������Q������R�   k���0�R� �Ѓ�������%�   t6������ u-��P����f4��P������Q�   k�	��0�Q� �Ѓ���������gu:������%�   u-��P���� 4��P������Q�   ����0�P� �Ѓ����������-u ������   ��������������������������R��������������  ��������@������ǅ����
   �   ǅ����
   �   ǅ����   ǅ����   �
ǅ����'   ǅ����   ��������   t2�   k� Ƅ����0��������Q�   �� ������ǅ����   �)ǅ����   ������%�   t��������   �������������� �  t�EP�������������������   ��������   t�UR�������������������   �������� tE��������@t�UR�B���������������������EP�&���������������������@��������@t�UR����������������������EP�������3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ������������������ }ǅ����   �%���������������������   ~
ǅ����   �����������u
ǅ����    �   i��  �������������������������������������������� �������������   �������RP������R������P�1�����0�������������RP������Q������R�m���������������������9~���������������������������������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0�������������������� �b  ��������@tv��������   t�   k� Ƅ����-ǅ����   �L��������t�   k� Ƅ����+ǅ����   �%��������t�   k� Ƅ���� ǅ����   ������+�����+�������`�����������u������Q�UR��`���Pj �
  ����p���Q������R�EP������Q������R�
  ����������t'��������u������R�EP��`���Qj0�+
  �������� ��   ������ ��   ǅ0���    ��������h�����������d�����d�����������d�������d��������� ��   ��h���f�f��z�����z���Rj�E�P��(���Q�|(������0�����h�������h�����0��� u	��(��� uǅ���������*��p���P������Q�UR��(���P�M�Q�	  ���N����(��p���R������P�MQ������R������P�c	  �������� |'��������t������R�EP��`���Qj ��  �������� tj������R�������ǅ����    �i��������� t������tǅ ���    �
ǅ ���   �� ������������� u&hh�h�Yj h�  hx�j��������u̃���� uF��%���    j h�  hx�h��hh��Q����ǅ����������P����|������������������������P����]����������M�3�������]Ë�\4�5�5l6�6�6.7�836D6"66X6g6 �I �7g8k7x8�8 ��<�8K:$?�9�<�8�>�;�??j:?0?�B   	
����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP������E��}��u�M�������U����M���]�������������������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��|�U�    �E�E��M���M�}� ~N�U��E��MQ�UR�E�P�w������M���M�U�:�u�E�8*u�MQ�URj?�L�������띋E�8 u�M�U���]������������������������������������������������U��Q�����9�u	�E�   ��E�    �E���]����������������������U��Q�E�E��M�Q�UR�EP�X�������]���������������U��Q�E�E��M�Qj �UR�f������]�����������������U��Q�E�E��M�Q�UR�EP�4������]���������������U��Q�E�E��M�Q�UR�EP��������]���������������U��������9�u	�E�   ��E�    �M��M�} t������U���E�    �E����E��]���������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h��h�Yj j6h��j�I�������u̃}� u.����    j j6h��h0�h������������   �U�U������    �� �Pj�������E�    �����    �� �P�K������EԋE�Pj �MQ����    �� �P�������E�����    �� �P�U�R������E������   ��a���    �� �Pj�;����ËE܋M�d�    Y_^[��]������������������������������������������������������������������������������������������������U��Q�E�E��M�Qj �UR� ������]�����������������U��� �E������EP�M��l����M����P�MQ�M������BtP�MQ�U�R�5�����E�}� u�E��E���E������M��M��M��d����E���]�������������������������������U���H�} u�} v�} t	�E�     3��  �} t	�M������}���w	�E�   ��E�    �U��U�}� u#h@�h�Yj jJhx�j��������u̃}� u0�����    j jJhx�h��h@��T�����   �  �MQ�M��4����M��z����   �����    �  �M���   ~C�} t�} v�URj �EP�:������r��� *   �g����M܍M������E��  �} ��   �} v	�E�   ��E�    �U��U�}� u#hvh�Yj j]hx�j��������u̃}� u=����� "   j j]hx�h��hv�U�����E�"   �M������E��}  �M�U��} t	�E�    �E�    �M��X����E��O  �B  �E�    �M�Qj �UR�EPj�MQj �M��*����BP� �E��}� t
�}� ��   �}� ��   �� ��z��   �} t�} v�MQj �UR�������3�t	�E�   ��E�    �M�M��}� u#h��h�Yj j{hx�j��������u̃}� u:����� "   j j{hx�h��h���!�����E�"   �M��R����E��L���� *   ���� �E̍M��0����E��*�} t�M�U���E�    �M������E���M�������]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�����j �EP�
��P�MQ�U�R�������E�}� u�E��E���E������E���]������������������������U��j �EP�MQ�UR�EP�L�����]�����������������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� �������������������������������������������U���$�E=��  u	f�E�)  �MQ�M������M�������   �����    u>�M��A|�U��Z�E�� �E���M�M�f�U�f�U��M��y���f�E���   �E=   }Yj�MQ�������uf�Uf�U��M��B���f�E��   �+�M��3��� �M���   f�
f�E��M�����f�E��`j�M�Qj�URh   �M������ �   �ዔ�   R��������uf�Ef�E��M������f�E��f�M�f�M�M�����f�E��]������������������������������������������������������������������������������������������U��j �EP������]�������������U��j
j �EP������]������������U��EPj
j �MQ�	����]��������U��EP�MQ� �����]������������U��EPj
j �MQ������]��������U��EPj
j �MQ�+	����]��������U��EP������]����������������U��j
j �EP�������]������������U��j
j �EP�4�����]������������U��j j j�EP�MQ�UR��
����]������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j�������E�    �EP�MQ�UR�EP�MQ�UR�[   ���E��E������   �j������ËE�M�d�    Y_^[��]����������������������������������������U����} t	�E�   ��E�    �E�E��}� u&h��h�Yj hX  h �j���������u̃}� u3�(���    j hX  h �h�h��������   �G  �U�    �} t	�E�     �} t	�E�   ��E�    �M�M�}� u&h0�h�Yj h^  h �j�N�������u̃}� u3����    j h^  h �h�h0��������   �   �EP�1������E��}� u3��   �M�Q���������E��UR�EP�MQj�U�R�;������M��U�: u����    ����� �Ej hr  h �h�hX��E�P�M�Q�U�P�����P�C������} t�M�U��3���]�������������������������������������������������������������������������������������������������������������������������������U���� ��E��=p� u3���   �}� u"�=� t�u����t3���   � ��M��}� ��   �} ��   �UR�������E��E��8 ��   �M��R������;E���   �E���U����=uo�M�Q�UR�E��Q���������uUh�  �U���M��TR�X����=�  r&h��h�Yj h�   h �j���������u̋M���E��D��M����M��O���3���]���������������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E�}� u&hl�h�Yj h�   h �j�'�������u̃}� u3�h���    j h�   h �h��hl��������   �%  �U�    �} t�} w�} u�} t	�E�    ��E�   �E��E�}� u&h��h�Yj h�   h �j��������u̃}� u3��
���    j h�   h �h��h���&�����   �   �} t�U� �EP�b������E��}� u3��d�M�Q�K��������U��} u3��F�E�;Mv�"   �5j h�   h �h��h���U�R�EP�MQ�Y����P������3���]�����������������������������������������������������������������������������������������������������������������U��j�h8�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} t	�E�   ��E�    �E�E��}� u#h��h�Yj jNh �j���������u̃}� u-�	���    j jNh �h��h���w����3���   h�  �UR�������=�  s	�E�   ��E�    �E܉E؃}� u#h��h�Yj jOh �j�O�������u̃}� u*����    j jOh �h��h���� ����3��<j�������E�    �UR�*������E��E������   �j�9�����ËEԋM�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������U��j�hX�h�Ld�    P���SVW���1E�3�P�E�d�    �E�    j�������E�    �EP�MQ�UR�EP�������E��E������   �j�<�����ËE�M�d�    Y_^[��]������������������������������������������������U���EP�MQ�������]����������U���EP�MQ������]����������U��Q�E=��  u3��G�M��   }�U���P�M#��&�U�Rj�EPj� ��u3�f�M��E��U#�]�����������������������������������U���$�} t�} v	�E�   ��E�    �E��E�}� u#hUh�Yj jh��j蔿������u̃}� u0�����    j jh��h�hU�2������   �-  �E�    �U�U�} tI�E���t?�U����U��E�;Er�  �M�Uf�f��M���M��:   �E�f��M���M�U�U��}� ��   �E������   �U����U��E�;Er��  �M�U�f�f��M���M�U����U��E����uU����U��E����/t5�U����\t*�M����M��U�;Ur�c  �\   �M�f��U���U�E�E��}� t@�M����t6�E����E��M�;Mr�#  �U�E�f�f�
�U���U�E����E����M�M��}� t�U����t5�M����.t*�E����E��M�;Mr��   �.   �E�f��M���M�U����t6�M����M��U�;Ur�   �E�M�f�f��E���E�M����M����U����U��E�;Ev�e3ɋU�f�
�}�tP�}���tG�E�;Es?�M+M�9h�s�h��U��	�E+E��E�M���Qh�   �U��E�PQ�$�����3���   3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R�������� L��t3�t	�E�   ��E�    �U��U܃}� u#hPLh�Yj jlh��j�i�������u̃}� u-���� "   j jlh��h�hPL�������"   ��   ��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���H�E�    �E�    �E�    �} u�e  �} u�} u�} t�} u�H  �} u�} u�} t�} u�+  �} u�}  u�} t�}  u�  �}$ u�}( u�}$ t�}( u��  �}� ��   �E�   �E�E��}� v�M����t�E���E�M����M��܋U����:u2�} t!�}s�  j�MQ�UR�EP��������M����M�_�} tY3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E�M���Qh�   �U��R��������E�    �E�    �E�E��	�M����M��U����t4�M����/t�E����\u�U����U���E����.u�U��U�빃}� t>�} t0�E�+E���E��M;M�w�  �U�R�EP�MQ�UR��������E��E�_�} tY3ɋUf�
�}�tK�}���tB�}v<�E��9h�s�h��M��	�U���U�E���Ph�   �M��Q��������}� ty�U�;Urq�} t0�E�+E���E��M ;M�w��   �U�R�EP�M Q�UR�,������}$ t0�E�+E����E��M(;M�w�   �U�R�E�P�M(Q�U$R��������   �} t0�E�+E���E��M ;M�w�   �U�R�EP�M Q�UR�������}$ tX3��M$f��}(�tJ�}(���tA�}(v;�U(��9h�s
�h��E��	�M(���M��U���Rh�   �E$��P�������3��  �E�   �} t_�} vY3ɋUf�
�}�tK�}���tB�}v<�E��9h�s�h��M��	�U���U܋E���Ph�   �M��Q�M������} t_�} vY3ҋEf��}�tK�}���tB�}v<�M��9h�s�h��U��	�E���E؋M���Qh�   �U��R��������} t^�}  vX3��Mf��} �tJ�} ���tA�} v;�U ��9h�s
�h��E��	�M ���MԋU���Rh�   �E��P�������}$ t_�}( vY3ɋU$f�
�}(�tK�}(���tB�}(v<�E(��9h�s�h��M��	�U(���UЋE���Ph�   �M$��Q�������} t	�E�   ��E�    �ỦUȃ}� u&h(�h�Yj h�   hX�j�ȵ������u̃}� u3�	����    j h�   hX�h��h(��c������   �   �}� t|3�t	�E�   ��E�    �U��U��}� u&h��h�Yj h�   hX�j�C�������u̃}� u0�����    j h�   hX�h��h����������   ��T���� "   �"   ��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��=,��t�=,��t�,�P�� ]��������������U��j j jj jh   @h(��T�,�]�������������U���<�E�    �E�    �E�H��pt	�U��pu'�E�H�U;�u	�E�   ��E�    �E��  �E�H��st�U�B��St	�E�    ��E�   �M��M��U��st�E��St	�E�    ��E�   �M�M��}� u�}� t[�U�;U�uD�E�H�� u	�E�   ��E�    �U�� u	�E�   ��E�    �E�;E�u	�E�   ��E�    �E���  �M�Q��dtv�E�H��itj�U�B��ot^�M�Q��utR�E�H��xtF�U�B��Xt:�M��dt1�U��it(�E��ot�M��ut�U��xt�E��X�,  �M�Q��dtE�E�H��it9�U�B��ot-�M�Q��ut!�E�H��xt�U�B��Xt	�E�    ��E�   �M��dt6�U��it-�E��ot$�M��ut�U��xt�E��Xt	�E�    ��E�   �M�;M�t3��   �U�B%   t	�E�   ��E�    �M��   t	�E�   ��E�    �U�;U�u;�E�H�� t	�E�   ��E�    �U�� t	�E�   ��E�    �E�;E�t3���M�;Uu	�E�   ��E�    �Eċ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE�ǅ ���    ǅ����    ǅ����    ǅ����    ǅ`���    ǅ���    ǅ8���    ǅ����    ǅP���    �EP��h���詸��ǅ����    ǅx���    ǅ����    ǅ����    ǅ��������ǅ��������ǅ��������ǅ��������ǅ��������ǅT���    ������������} tǅ���   �
ǅ���    ����������������� u&h �h�Yj h  hx�j�#�������u̃����� uI�a����    j h  hx�h<�h �������ǅ����������h����������������6  �} tǅ����   �
ǅ����    ������������������ u&h��h�Yj h  hx�j�z�������u̃����� uI�����    j h  hx�h<�h��������ǅ���������h����=���������16  ǅ����    �U������ǅ����    �����������������������5  ������u������ u��5  ǅ����    ǅd���    ǅT���    ǅ ���    ǅ��������ǅ����    ǅ����    �������Mǅ��������ǅ��������ǅ��������ǅ���������Uf�f������������������U���U����� �N2  ������ �A2  �������� |%��������x��������(����������
ǅ����    ������������k�����	��d�����H�����d�����d�����  �U���%��  �������u\j
��x���Q�UR�B�������~9��x������$u+������ uh@  j ������R�a�����ǅ����   �
ǅ����    �������.  j
��x���P�MQ�����������������x������U������ ��   ������ |#��x������$u������d}ǅ ���   �
ǅ ���    �� ��������������� u&h�h�Yj hU  hx�j自������u̃����� uI������    j hU  hx�h<�h�������ǅ����������h����J����������>3  ������;�����~�����������������������������������   ��d�����   3�tǅ����   �
ǅ����    ���������������� u&h��h�Yj ha  hx�j蚩������u̃���� uI������    j ha  hx�h<�h���2�����ǅ����������h����]����������Q2  ��d����������������I/  �������$��������� u	������t������u�������u�/  ǅP���   ������Q�UR������P�A  ����.  ǅ���    �������8�����8�����������������`���ǅ����    ǅ��������ǅP���    �.  ������������������ ����������wj���������$�̮���������������E���������������4���������������#�������ʀ   ����������������������.  ��������*��  ������ u�UR虾�����������  j
��x���P�MQ�d���������������x������U������ �)  ������ |#��x������$u������d}ǅ���   �
ǅ���    ����������������� u&h �h�Yj h�  hx�j��������u̃����� uI�P����    j h�  hx�h<�h �������ǅ���������h���������������/  ������;�����~�������� ������������ ����� ����������������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R�)�������tǅ����   �
ǅ����    ������������������ u&h��h�Yj h�  hx�j賥������u̃����� uI������    j h�  hx�h<�h���K�����ǅ����������h����v����������j.  �v+  �+����������������H�����H���Q�	����������������� }���������������������؉������k�����
�������DЉ������+  ǅ����    ��*  ��������*��  ������ u�UR芻�����������  j
��x���P�MQ�U���������������x������U������ �)  ������ |#��x������$u������d}ǅ����   �
ǅ����    ������������������ u&h��h�Yj h�  hx�j��������u̃����� uI�A����    j h�  hx�h<�h��������ǅ����������h����ƽ���������,  ������;�����~��������������������������������������������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R��������tǅ<���   �
ǅ<���    ��<��������������� u&h8�h�Yj h�  hx�j褢������u̃����� uI������    j h�  hx�h<�h8��<�����ǅ ���������h����g����� ����[+  �g(  �+��������������������������Q������������������� }
ǅ���������k�����
�������LЉ������(  ��������(�����(�����I��(�����(���.�D  ��(�������$����E���lu�U���U������   �����������������������   �U���6u,�M�Q��4u �E���E�������� �  �������   �U���3u)�M�Q��2u�E���E������������������e�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu��������   �������ǅd���    �����#�������� ���������������   �������&  ��������0�����0�����A��0�����0���7��#  ��0�����x��$�<�������%0  u�������� ������ǅP���   ������ u�UR�ض����f��|����   ������ |������d}ǅ����   �
ǅ����    ������������������ u&h��h�Yj hz  hx�j蕟������u̃����� uI������    j hz  hx�h<�h���-�����ǅ@���������h����X�����@����L(  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R���������tǅ4���   �
ǅ4���    ��4��������������� u&h��h�Yj h~  hx�j�]�������u̃����� uI�����    j h~  hx�h<�h���������ǅ����������h���� ����������'  �w!  �,������������������������Q賴����f��|����������� ��   ��|���%�   �   k� ��@���ǅ����   ������s��`���������Ƅ@��� ��h�������P��h����}�����QtR��@���P������Q�|�������}
ǅ8���   ��   k� f��|���f������������������ǅ����   �   ������ u�EP�г������L����  ������ |������d}ǅ����   �
ǅ����    ��������,�����,��� u&h��h�Yj h�  hx�j莜������u̃�,��� uI������    j h�  hx�h<�h���&�����ǅ����������h����Q����������E%  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������P������Qj��������������P���������tǅ����   �
ǅ����    ������������������ u&h��h�Yj h�  hx�j�V�������u̃����� uI�����    j h�  hx�h<�h���������ǅ8���������h���������8����$  �p  �+��������������������������R謱������L�����L��� t��L����x u#�p�������������R��������������d������%   t/��L����Q��������L���� �+���������ǅP���   �(ǅP���    ��L����Q��������L�����������  ��������0  u�������� �������������uǅ����������������������������,��������� u�EP覰�����������  ������ |������d}ǅ$���   �
ǅ$���    ��$��������������� u&h��h�Yj h:  hx�j�d�������u̃����� uI�����    j h:  hx�h<�h���������ǅ����������h����'����������"  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������P������Qj��������������P��������tǅ����   �
ǅ����    ��������|�����|��� u&h��h�Yj h>  hx�j�,�������u̃�|��� uI�j����    j h>  hx�h<�h���������ǅ����������h���������������   �F  �+����������������0�����0���R肮������������������ ��   ������ u�p���������������H���ǅ����    ���������������������;�,���}O��H������tB��h����E���P��H����R�R�������t��H�������H�����H�������H�����   ������ u�t�������ǅP���   ��������$�����,�����x�����,�������,�����x��� t��$������t��$�������$���뾋�$���+���������������  ������ u�MQ�4�����������  ������ |������d}ǅ���   �
ǅ���    �������t�����t��� u&h��h�Yj h�  hx�j��������u̃�t��� uI�0����    j h�  hx�h<�h��������ǅ���������h���赯��������  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������Q������Rj��������������Q�0�������tǅ����   �
ǅ����    ��������l�����l��� u&h��h�Yj h�  hx�j躔������u̃�l��� uI������    j h�  hx�h<�h���R�����ǅp���������h����}�����p����q  ��  �+����������������(�����(���P��������������������   3�tǅ���   �
ǅ���    �������d�����d��� u&h�h�Yj h�  hx�j�ԓ������u̃�d��� uI�����    j h�  hx�h<�h��l�����ǅh���������h���藭����h����  ��  �������� t�����f������f��������������ǅ8���   �  ǅ���   �������� f��������������@��������������  ������ ��  ������ |������d}ǅ����   �
ǅ����    ��������\�����\��� u&h��h�Yj h�  hx�j蜒������u̃�\��� uI������    j h�  hx�h<�h���4�����ǅ����������h����_����������S  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������Q������Rj��������������Q���������tǅ���   �
ǅ���    �������T�����T��� u&h(�h�Yj h�  hx�j�q�������u̃�T��� uI�����    j h�  hx�h<�h(��	�����ǅ`���������h����4�����`����(  �  ������������ǅ ���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Yh�  hp�j������]  P訌������T�����T��� t ��T�����������������]  �� ����
ǅ�����   ������ u#�E���E�M�Q��A��������������!  ������ |������d}ǅ����   �
ǅ����    ��������L�����L��� u&h��h�Yj h  hx�j�ď������u̃�L��� uI�����    j h  hx�h<�h���\�����ǅ ���������h���臩���� ����{  ������t&h��h�Yj h  hx�j�C�������u̋������������������������������������Q��A���������������h����	���P�����Q������R������P�� ���Q������R������P�   k���0�P� �Ѓ���������   t6������ u-��h�������P������R�   k�	��0�R� �Ѓ���������gu;��������   u-��h����Z���P������R�   ����0�Q� �Ѓ����������-u!��������   ��������������������������P�������������R  ��������@������ǅD���
   �   ǅD���
   �   ǅ����   ǅ ���   �
ǅ ���'   ǅD���   ��������   t8�   k� �0   f��<����� �����Q�   �� f��<���ǅ`���   �)ǅD���   ��������   t������   �������������� �  �P  ������ u�UR�������������������%  ������ |������d}ǅ����   �
ǅ����    ��������D�����D��� u&h��h�Yj h�  hx�j�~�������u̃�D��� uI�����    j h�  hx�h<�h��������ǅX���������h����A�����X����5  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R輾������tǅ����   �
ǅ����    ������������������ u&h�h�Yj h�  hx�j�F�������u̃����� uI�����    j h�  hx�h<�h��������ǅ���������h����	����������  �`  �1����������������P�����P���Q��������������������  ��������   �P  ������ u�EP谹�����������������%  ������ |������d}ǅ����   �
ǅ����    ������������������ u&h��h�Yj h�  hx�j��������u̃����� uI�Z����    j h�  hx�h<�h��������ǅ���������h����ߣ���������  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������P������Qj��������������P�Z�������tǅ����   �
ǅ����    ������������������ u&h��h�Yj h�  hx�j��������u̃����� uI�"����    j h�  hx�h<�h���|�����ǅ����������h���觢���������  ��  �1��������������������������R膷�����������������z	  �������� ��  ��������@�T  ������ u�UR����������������������'  ������ |������d}ǅ����   �
ǅ����    ������������������ u&h��h�Yj h�  hx�j謇������u̃����� uI������    j h�  hx�h<�h���D�����ǅ����������h����o����������c  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R��������tǅ����   �
ǅ����    ������������������ u&h��h�Yj h�  hx�j�t�������u̃����� uI�����    j h�  hx�h<�h��������ǅ����������h����7����������+  �	  �3��������������������������Q�ʜ�������������������S  ������ u!�UR袜��������������������)  ������ |������d}ǅx���   �
ǅx���    ��x�����p�����p��� u&h��h�Yj h�  hx�j�V�������u̃�p��� uI�����    j h�  hx�h<�h���������ǅ����������h��������������  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������R������Pj��������������R蔷������tǅh���   �
ǅh���    ��h�����`�����`��� u&h��h�Yj h  hx�j��������u̃�`��� uI�\����    j h  hx�h<�h��������ǅ����������h���������������  �8  �5����������������|�����|���Q�t���������������������  ��������@�R  ������ u�EP�;�������������������&  ������ |������d}ǅX���   �
ǅX���    ��X�����P�����P��� u&h��h�Yj h  hx�j��������u̃�P��� uI�0����    j h  hx�h<�h��������ǅt���������h���赜����t����  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������P������Qj��������������P�0�������tǅH���   �
ǅH���    ��H�����@�����@��� u&h��h�Yj h  hx�j躁������u̃�@��� uI������    j h  hx�h<�h���R�����ǅl���������h����}�����l����q
  ��  �2����������������d�����d���R��������������������O  ������ u�EP������3ɉ������������'  ������ |������d}ǅ8���   �
ǅ8���    ��8�����0�����0��� u&h��h�Yj h4  hx�j蟀������u̃�0��� uI������    j h4  hx�h<�h���7�����ǅ\���������h����b�����\����V	  ������ �2  �������������� uG��������Ǆ����   ��������f������f����������������������������   ������Q������Rj��������������Q�ݲ������tǅ(���   �
ǅ(���    ��(��������������� u&h��h�Yj h8  hx�j�g������u̃����� uI�����    j h8  hx�h<�h���������ǅT���������h����*�����T����  �  �3����������������L�����L���P轕����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�X�����\�����������   ���������������X�����������\����������� �  u(������%   u��X�����\����� ��X�����\��������� }ǅ����   �%���������������������   ~
ǅ����   ��X����\���u
ǅ`���    �   i��  ��������������������D�������������������D��� ��X����\�����   ��D����RP��\���R��X���P������0��4�����D����RP��\���Q��X���R�H�����X�����\�����4���9~��4���� �����4�����������4�������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0��������������������u������ u�  ��8��� �a  ��������@��   ��������   t!�   k� �-   f��<���ǅ`���   �V��������t!�   k� �+   f��<���ǅ`���   �*��������t�   k� �    f��<���ǅ`���   ������+�����+�`�����������������u������Q�UR������Pj ��  ��������Q������R�EP��`���Q��<���R��  ����������t'��������u������R�EP������Qj0�l  ����P��� ��   ������ ��   �����������������������������<�����������������<��� ��   ��h��������P��h��������� �HtQ�����R��|���P�ھ���������������� ǅ���������2������Q�UR��|���P�)  ������������������X����(������R������P�MQ������R������P�  �������� |'��������t������R�EP������Qj �8  ����T��� tj��T���R苈����ǅT���    ������d��� t��d���tǅ����    �
ǅ����   ������������������ u&hh�h�Yj h�  hx�j�~y������u̃����� uI輿���    j h�  hx�h<�hh�������ǅ4���������h����A�����4����5  �������  ������ ��  ǅ����    ���������������������;�������  ��������������������������������������   ������$������������E�������MQ�[������d  ���������E�������MQ�7������@  ���������E�������MQ�_������  ���������E�������MQ�;�������   ���������E�������MQ�ˎ������   ���������E�������MQ��������������������   3�tǅ����   �
ǅ����    ������������������ u&h��h�Yj h2	  hx�j�mw������u̃����� uF諽���    j h2	  hx�h<�h��������ǅ,���������h����0�����,����'����������������$�����h���������$����M�3�豕����]�s|�|}�}�������r}�}a}P}�}�} �I ����� �R�V�d����m�r��� �S����җ���   	
��7�[��ӭ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E�H��@t�U�z u�E����U�
�4�EP�MQ舦�����Ё���  u�E� ������M����E�]�������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�U������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��~�U�    �E�E��M���M�}� ~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������뛋E�8 u�M�U���]����������������������������������������������U���  ���3ŉE�ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    �EP��d�����n��ǅ����    �f�����P����} tǅ0���   �
ǅ0���    ��0�����`�����`��� u&h �h�Yj h  hx�j�d������u̃�`��� uI������    j h  hx�h\�h ��U�����ǅ���������d����~��������  �} tǅ(���   �
ǅ(���    ��(����� ����� ��� u&h��h�Yj h  hx�j�d������u̃� ��� uI�R����    j h  hx�h\�h��謢����ǅ���������d�����}���������  ǅ����    ǅ����    ǅ����    ǅ����    ǅt���    �Uf�f������������������U���U����� ��  ������ ��  �������� |%��������x��������(�����<����
ǅ<���    ��<���������k�����	��������H�����������������   3�tǅ8���   �
ǅ8���    ��8�����T�����T��� u&h��h�Yj he  hx�j�b������u̃�T��� uI�ʨ���    j he  hx�h\�h���$�����ǅ����������d����O|���������n  ��������,�����,�����  ��,����$���ǅ����   ������Q�UR������P�  ���J  ǅ����    ������������������������������������ǅ����    ǅ��������ǅ����    ��  �������������������� ������������wj����������$������������������E���������������4���������������#�������ʀ   ����������������������e  ��������*u:�UR��w���������������� }���������������������ى������k�����
�������LЉ������  ǅ����    ��  ��������*u'�EP�Ow���������������� }
ǅ���������k�����
�������DЉ������  ��������������������I������������.�1  ��������8��$�$��U���lu�M���M��������   �����������������������   �M���6u+�E�H��4u�U���U������ �  �������   �M���3u(�E�H��2u�U���U������%����������S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    ������#�������� ���������������   �������D  ��������������������A������������7��
  �����������$�h���������0  u�������� ������ǅ����   �EP�Hu����f�������������� ��   ���������   �   k� ������ǅL���   ��L���s��������L���Ƅ���� ��d�������P��d�������� �HtQ������R������P��������}
ǅ����   ��   k� f������f������������������ǅ����   �s	  �UR�mt���������������� t�������x u#�p�������������R荇�����������d������%   t/�������Q������������� �+���������ǅ����   �(ǅ����    �������Q���������������������  ��������0  u�������� �������������uǅ4���������������4�����4����������EP�ps������������������ ��   ������ u�p�������������������ǅ����    ���������������������;�����}O���������tB��d����3���P�������P�@�������t������������������������������   ������ u�t�������ǅ����   ������������������������������������������ t���������t��������������뾋�����+��������������2  �UR�,r������\�����������   3�tǅD���   �
ǅD���    ��D�����$�����$��� u&h�h�Yj h�  hx�j��Z������u̃�$��� uI�.����    j h�  hx�h\�h�舙����ǅ ���������d����t���� �����	  �g  �������� t��\���f������f����\����������ǅ����   �-  ǅ����   �������� f��������������@������������������ǅt���   ������ }ǅ����   �7������ u��������guǅ����   �������   ~
ǅ����   �������   ~Yh�  hp�j������]  P��U���������������� t ��������������������]  ��t����
ǅ�����   �E���E�M�Q��A���������������d����S���P������Q������R������P��t���Q������R������P�   k���0�P� �Ѓ���������   t6������ u-��d�������P������R�   k�	��0�R� �Ѓ���������gu;��������   u-��d���褥��P������R�   ����0�Q� �Ѓ����������-u!��������   ��������������������������P�`�������������  ��������@������ǅ����
   �   ǅ����
   �   ǅ����   ǅ����   �
ǅ����'   ǅ����   ��������   t8�   k� �0   f��������������Q�   �� f������ǅ����   �)ǅ����   ��������   t������   �������������� �  t�UR�i������������������   ������%   t�MQ�?������������������   �������� tE��������@t�MQ��m��������������������UR�m��������������������@��������@t�MQ�{m�������������������UR�`m����3ɉ�������������������@tG������ >|	������ s3�������؋������� �ى�������������������   ��������������������������������������� �  u(������%   u�������������� ������������������ }ǅ����   �%���������������������   ~
ǅ����   �����������u
ǅ����    �   i��  ������������������������������������������ �������������   �������RP������R������P�n����0�������������RP������Q������R��l��������������������9~���������������������������������������������@����   i��  ������+���������������������������������   tG������ t�   k� �������
��0t'���������������������0�������������������� �a  ��������@��   ��������   t!�   k� �-   f������ǅ����   �V��������t!�   k� �+   f������ǅ����   �*��������t�   k� �    f������ǅ����   ������+�����+�������x�����������u������Q�UR��x���Pj �	  ����P���Q������R�EP������Q������R��	  ����������t'��������u������R�EP��x���Qj0�F	  �������� ��   ������ ��   ��������|����������������������������������������������� ��   ��d���衟��P��d���蕟��� �HtQ��|���R������P蔖������X�����X��� ǅ���������2������Q�UR������P�  ����|����X�����|����X����(��P���R������P�MQ������R������P�  �������� |'��������t������R�EP��x���Qj �  �������� tj������R�E`����ǅ����    ���������� t������tǅH���    �
ǅH���   ��H�����@�����@��� u&hh�h�Yj h�  hx�j�8Q������u̃�@��� uF�v����    j h�  hx�h\�hh��Џ����ǅ���������d�����j���������������������d�����j��������M�3��o����]Ð�����������R���W�h�F�5�|��� �I ���������� �6���������Q��j�1�	���������c�   	
��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��E�H��@t�U�z u�E����U�
�4�EP�MQ�h������Ё���  u�E� ������M����E�]�������������������������������������U��Q�E�E��M���M�}� ~!�UR�EP�MQ�U������U�:�u��ʋ�]�������������������U����E��M�U�B��@t�M�y u�U�E�M��~�U�    �E�E��M���M�}� ~P�Uf�f�E��MQ�UR�E�P��������M���M�U�:�u�E�8*u�MQ�URj?��������뛋E�8 u�M�U���]����������������������������������������������U���4���3ŉE�V�E�H��@�d  �UR��{�������t@�EP�{�������t/�MQ�{���������UR�{���������0��E���E���E��H$�����у�tj�EP�`{�������t@�MQ�O{�������t/�UR�>{���������EP�-{���������0��E���E���MԊQ$������uh�M�Q���U�E�M�H�}� |2�U�f�Mf��U����  f�U�E����U�
f�E��  ��EP�MQ�k�����  �(  �UR�z�������t@�EP�}z�������t/�MQ�lz���������UR�[z���������0��E���E���E��H��   ��   �URj�E�P�M�Q�'�������t
���  ��   �E�    �	�U����U��E�;E�}s�M�Q���U؋E�M؉H�}� |.�U��M��T��E�����   �U�E����U�
��EP�M��T�R�h������E�}��u���  �k�|����E%��  �[�E�H���M܋U�E܉B�}� |/�M�f�Ef��M����  f�M�U����M�f�E����UR�EP�j����^�M�3��_d����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�hx�h�Ld�    P���SVW���1E�3�P�E�d�    3�f�E�} t	�E�   ��E�    �M܉M؃}� u#h��h�Yj j3h��j�ZD������u̃}� u-蛊���    j j3h��h��h������������  �M�E�E��M�Q�ez�����E�    �U�R�EP�g�����f�E��E������   ��M�Q�������f�E�M�d�    Y_^[��]��������������������������������������������������������������������U��EP�MQ�i����]�����������U����E�E�M�M��E�    �	�U����U��}�}�E��M���E����E��M���M��Ӌ�]���������������������U��Q�E�    �	�E����E��}�}�M��U��    ���]������������������U����E�������E��E%  �yH���@�   +ȉM��   �M���U��E��M��R�E�P�M��U��P��K�����E��M����M��	�U����U��}� |)�}� t#�E��M��Rj�E��M��R�K�����E��ȋE���]���������������������������������������������������������U��Q�E�    �	�E����E��}�}�M��U�<� t3���߸   ��]��������������������������U����E�    �E���E��M����M�E��������E��U��  �yJ���B�   +E�   �M���U�E��M��#U�t'�E�P�MQ�*o������u�U�R�EP��m�����E����M���E��M#��E��M���U����U��	�E����E��}�}�M��U��    ��E��]�������������������������������������������������������������U���V�E�������E��E%  �yH���@�E�����M����҉U��E�    �E�    �	�E����E��}�}M�M��U��#E�E�M��U���M���M��U���E��M��U�E��M���    +M��U���U���E�   �	�E����E��}� |.�M�;M�|�U�+U��E��M�u������E��M��    ��^��]���������������������������������������������������������������������U����E�������E��E%  �yH���@�   +ȉM�����M����҉U�E��M��#U�t3��1�E����E��	�M����M��}�}�U��E�<� t3���߸   ��]�����������������������������������������������U����E�    �EE�E��M�;Mr�U�;Us	�E����E��M�U���E���]�������������������U���@���3ŉE��E�H
���  ���?  �M��U�B
% �  �E��   k� �E�H�L�   �� �E�H�L��U����   ��D��}����u8�E�    �U�R��W������t	�E�    ��E�P�[�����E�   �  �M�Q�U�R�S������E��E̋M�QR�E�P�zw������t	�M����M��U�E�J+H9M�}�U�R�:[�����E�    �E�   �  �E�M�;Hn�U�R�E�P�������M̉M��U�B+E��EȋM�Q�U�R�ly�����E�HQ�U�R��v�����E�H��Q�U�R�Cy�����E�    �E�   �   �E�M�;|T�U�R�Z�����   k� �T���   ��   k� �T��U�BP�M�Q��x�����U��MA�E��E�   �C�U�E�B�Eع   k� �D�%����   k� �D��E�HQ�U�R�x�����E�    �E�H���    +щUă}� t	�E�   ���E�    �   k� �E؋M���D�EԉEЋM�y@u�U�EЉB�   �� �U�D����M�y u�U�EЉ�E܋M�3��eZ����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��h0��EP�MQ�������]�������U��hH��EP�MQ�݁����]�������U������3ŉE��E�    �E�H
���  f�M�U�B
% �  f�E�   k� �E�H�L�   �� �E�H�L��U����   ��D�j@�U�R�#t������t�   k� �D�   �f�U�f��f�U��E�=�  u�E�   �   k� �E�L��H�   �� �E�L���U��E�ЋMf�Q�E�M�3��xX����]����������������������������������������������������������������������������U������3ŉE��EPj j j �MQ�UR�EP�M�Q�vw���� �E�UR�E�P�Or�����E�}�u	�M���M�E�M�3���W����]�����������������������������������������U���T���3ŉE�3�f�E��E�    �E�    �E�    �E�    �Mf�Q
f�U�Ef�H
f�M��U��E�3Ё� �  f�U��M���  f�M��U���  f�U��E��M��f�E��U���  }�E�=�  }�M����  ~9�U���t	�E� �����E� ���E�M��H�U�B    �E�     �  �M���?  "�U�B    �E�@    �M�    ��  �U��u9f�E�f��f�E�M�Q�����u�E�x u�M�9 u3ҋEf�P
�  �M��uMf�U�f��f�U�E�H�����u3�U�z u*�E�8 u"�M�A    �U�B    �E�     �R  �E�    �E�    �	�M؃��M؃}���   �U���U��E�   �   +E؉E��	�Mȃ��Mȃ}� ~x�UỦU��EEԉE��M܍T��U��E���U���ȉM��M�Q�U�R�E��Q��?�����E��}� t�U�f�D�f���M�f�D�Ũ��ŰEԃ��E��y����M܃��M��<����U���?  f�U��E��~%�M���   �u�U�R�<����f�E�f��f�E����M��Qf�U�f��f�U��E��},�M���t	�UЃ��UЍE�P�O5����f�M�f��f�M��̃}� t�U���f�U��E�= �  �M����� �� � u_�}��uP�E�    �}��u8�E�    �U�����  u� �  f�E�f�M�f��f�M��f�U�f��f�U��	�E����E��	�M���M��U���  |6�E���t	�E� �����E� ���M�UĉQ�E�@    �M�    �-�Uf�E�f��M�U�Q�E�M��H�U��E�ЋMf�Q
�M�3��S����]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U������3ŉE��p���`�E�} u�   �} }�M�ىM�и��`�U�} u3��Mf��} tp�U��T�U�E���E�M���M�}� u��kU�U�U�E���� �  |#�U��E��J�M�R�U��E���E�M��M�U�R�EP��t����늋M�3��Q����]����������������������������������������������������������������U����E���   �t	�E�   ��E�    �U��U�E�H��   �t	�E�   ��E�    �U��U��E���U�
�E�H��M�U�J�E�H��M��U�J��]����������������������������������U����E�H��t	�E�   ���E�    �U��U�E�H��t	�E�   ���E�    �U��U��E�H��U�J�E�H��M�U�J�E���M��U�
��]���������������������������������������U���   ���3ŉE��E��E�3�f�M�ǅl���   �E�    �E�    �E�    ǅp���    �E�    ǅ|���    �E�    �E�    �E�    �E�    3�f�U�3�f�E��E�    �E�    �}$ tǅh���   �
ǅh���    ��h�����\�����\��� u#h��h�Yj j~h�j�0������u̃�\��� u-��v���    j j~h�h��h���-o����3��  �E�E̋M̉M��	�Ũ��ŰE���� t!�U����	t�M����
t�E����u�Ƀ}�
�;  �Ů�EӋM̃��M̋Uȉ�`�����`����  ��`����$����MӃ�1|�UӃ�9�E�   �Ẽ��E��   �MӋU$����   ��;�u	�E�   �`�Eӈ�t�����t���+t��t���-t#��t���0t�*�E�   �1�E�   3�f�M��"�E�   � �  f�U���E�
   �Ẽ��E��U  �E�   �MӃ�1|�UӃ�9�E�   �Ẽ��E��|�MӋU$����   ��;�u	�E�   �[�EӉE��M���+�M��}�:w5�U���8��$�(��E�   �+�E�   �"�M̃��M��E�   ��E�
   �Ũ��U��  �EӃ�1|�MӃ�9�E�   �Ũ��U��K�EӋM$����   ��
;�u	�E�   �*�Uӈ�T�����T���0t�	�E�   ��E�
   �E��E��5  �E�   ��M̊�UӋẼ��E��MӃ�0|:�UӃ�91�}�s �E����E��MӃ�0�U��
�E����E��	�M����M���UӋE$����   ��;�u	�E�   �R�MӉM��U���+�U��}�:w,�E������$�t��E�   �"�Ũ��U��E�   ��E�
   �Ẽ��E��`  �E�   �E�   �}� u'��M̊�UӋẼ��E��MӃ�0u�U����U�����E̊�MӋŨ��U��EӃ�0|8�MӃ�9/�}�s'�U����U��EӃ�0�M���U����U��E����E���MӉM��U���+�U��}�:w,�E������$����E�   �"�Ũ��U��E�   ��E�
   �Ẽ��E��z  �E�   �MӃ�0|�UӃ�9�E�   �Ẽ��E���E�
   �M��M��=  �Ũ��U��EӃ�1|�MӃ�9�E�	   �Ũ��U��X�Eӈ�x�����x���+t0��x���-t��x���0t�%�E�   �)�E�   ǅl���������E�   ��E�
   �M��M��  ǅp���   ��Ů�EӋM̃��M��UӃ�0u���EӃ�1|�MӃ�9�E�	   �Ũ��U���E�
   �Ẽ��E��R  �MӃ�1|�UӃ�9�E�	   �Ẽ��E��*�Mӈ�X�����X���0t�	�E�   ��E�
   �U��U���   ǅp���   �E�    ��E̊�MӋŨ��U��EӃ�0|,�MӃ�9#kU�
�EӍLЉM��}�P  ~	�E�Q  �뺋U��U���E̊�MӋŨ��U��EӃ�0|�MӃ�9���E�
   �Ũ��U��g�}  tQ�Ẽ��E��Mӈ�d�����d���+t��d���-t��E�   ǅl���������E�   ��E�
   �U��U���E�
   �Ẽ��E������M�Ủ�}� �`  �}� �V  ��|��� �I  �}�vF�   k��T���|�   k��T����   k��T��E�   �U����U��E����E��}� ��   �M����M��	�U����U��E����u�U����U��E����E��ٍM�Q�U�R�E�P�X������l��� }�M��ىM��U�U��U���p��� u	�E�E�E��}� u	�M�+M�M��}�P  ~	�E�   �E�}�����}ǅ|���   �0�UR�E�P�M�Q�^����f�U�f�U��E։E��MډM�f�U�f�U��3�f�E�3�f�M��UĉU��E��E��}� u$3�f�M�3�f�U��EĉE��M��M��U����U��Y�}� t(��  f�E��E�   ��E�    3�f�M��U����U��+��|��� t"3�f�E�3�f�M��UĉU��E��E��M����M��Uf�E�f��M�U��Q�E�M��H�U��E�ЋMf�Q
�E��M�3��gF����]Ë���i����^�D���l������W������� �  �7�.�I�  ���/�  �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   ���3ŉE��M  f�E��M   f�M���   f�U��E��C�E���E���E���E���E���E���E���E���E���E���E���E�?�E�   f�Ef�EЋM�M��U�U��E�% �  f�E��MЁ��  f�M��U̅�t	�E�@-��M�A �UЅ�uj�}� ud�}� u^3��Mf��Ú� �  u	�E�-   ��E�    �E�M��H�U�B�   k� �U�D
0�   �� �M�D �   ��  �UЁ��  �b  �   �Mf��}�   �u�}� tP�U���   @uEj jvh��h�h0�h��j�E��P��i����P�-�����M�A�E�    ��   �U̅�tT�}�   �uK�}� uEj j|h��h�h��h��j�E��P�{i����P�,�����M�A�E�    �   �}�   �uK�}� uEj h�   h��h�h��hD�j�U��R�$i����P�b,�����E�@�E�    �Cj h�   h��h�hP�h��j�M��Q��h����P�,�����U�B�E�    �\  �E���f�E��MЁ��   f��|����U���f�U��E��M����U��M�����U��M����+E��E��U���f�U�f�E�f�E��M��M��U��U�3�f�E�j�M���Q�U�R�V�����E�=�?  |f�M�f��f�MȍU�R�E�P�^b�����Mf�U�f��E��tn�M�M�M�} ^3ҋEf��Ḿ� �  u	�E�-   ��E�    �U�E��B�M�A�   k� �M�D0�   �� �E�D �   �.  �}~�E   �M����?  �M�3�f�U��E�    �	�E����E��}�}�M�Q�:&������}� }-�U��ځ��   �U��	�E����E��}� ~�M�Q��������U���UԋE���E��	�M����M��}� ~a�U��U؋E�E܋M��M��U�R��%�����E�P�%�����M�Q�U�R������E�P�%�����M���0�UԈ
�Eԃ��E��E� 됋Mԃ��MԋUԊ�EǋMԃ��M��Uǃ�5|_�	�Eԃ��EԋM��9M�r�U����9u�M��0�ًU��9U�s�Eԃ��EԋMf�f���Ef��MԊ���EԈ�   �	�Mԃ��MԋU��9U�r�E����0u�ߋU��9U�s[3��Mf��Ú� �  u	�E�-   ��E�    �E�M��H�U�B�   k� �U�D
0�   �� �M�D �   �&�U���E�+��M�A�U�B�M�D �E��M�3��<����]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����EP�M�R�E�Q�%�����E��}� t0�U��Rj�E�HQ�e%�����E��}� t�U�B���M�A�U��R�E�HQ�U�BP�0%�����E�}� t�M�Q���E�P�M��Q�U�BP�M�QR��$������]����������������������������������������������������U����E�    �E%�   t	�M����M��U��   t	�E����E��M��   t	�U����U��E%   t	�M����M��U��   t	�E����E��M��   t�U���   �U��E% `  �E��}� @  w�}� @  t$�}� t�}�    t#�:�}� `  t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��@�  �U�}�@t!�}� �  t&�}�@�  t�'�E�   �E���M���   �M���U���   �U��E���]�����������������������������������������������������������������������������������������������U��Q�E�    �E��?th�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]�����������������������������������������������U��Q�]��e���U��E�P�7�������]�����������������U����} t^��}��E�P�F  ���E��M#M�U��#U�ʉM�E�;E�t'�M�Q�,  ��f�E��m���}��U�R�  ���E�E�M��} t)�= �|�UR�EP�J   ���M��	�U�    �   ��]�����������������������������������������������U����E%�E�]��M�Q�������E��U#U�E��#E�ЉU�M�;M�u�E��+�U�R�s   ���E��E�P�������]��M�Q�D�������]������������������������������U��Q�E��  �E�P�������]����������������������U����E�    �E��t�M��ɀ   �M��U��t�E�   �E��M��t�U���   �U��E��t�M���   �M��U��t�E�   �E��M��   t�U���   �U��E%   �E��}�   w�}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U��� @  �U���E�    �E���M��� `  �M��U��   �U�}�   t�}�   t�}�   t�$�E�@�  �E���M���@�M���U��� �  �U��E���]�����������������������������������������������������������������������������������������������U��Q��<���E��E�P���������]���������������������U����E�    �E��t	�M����M��U��t	�E����E��M��t	�U����U��E��t	�M����M��U�� t	�E����E��M��t�U���   �U��E%   �E��}�   �}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��   �U�t*�}�   t�}�   t�"�E��E���M���   �M���U���   �U��E%   t�M���   �M��E���]�����������������������������������������������������������������������������������������U��Q�E�    �E��?tn�M��t	�U����U��E��t	�M����M��U��t	�E����E��M��t	�U����U��E�� t	�M����M��U��t�E�   �E��E���]����������������������������������������U��QV�}���= �|�E�P�3����������������M�Q������^��]������������������U�����}��E�P�L������E�M#M�U��#U�ʉM�E�;E�t'�M�Q�2  ��f�E��m���}��U�R�
������E�= �|B�EP�MQ�^������E��U�#���E�#��;�t�E�E�   ����E�E����E��]���������������������������������������������������U��E%����P�MQ�q7����]�������U����:��� �E�����Y���D����}� t/�M��Q�%  t �M��Q���U��E��@    �M��A��  ��]����������������������������U���3�f�E��M��t�U���f�U��E��t�M���f�M��U��t�E���f�E��M��t�U���f�U��E��t�M��� f�M��U��   t�E���f�E��M��   �M��}�   w�}�   t&�}� t�}�   t&�B�}�   t+�7f�U�f�U��-�E�   f�E���M���   f�M���U���   f�U��E%   �E�t�}�   t�}�   t"�(�M���   f�M���U���   f�U��f�E�f�E��M��   t�U���   f�U�f�E���]�����������������������������������������������������������������������������������������������������U����} 	 u>�}�u8��}��E�%=  ==  u$�= �|�]��M�����  ���  u�;��7j hN  h��h�h@��U������R�EPj � ����P��������]�����������������������������������������U�����}��E�P�������E��= �|�]�M�Q������E���E���]������������������U��Q�} t��}��E�P�������M��} t
������U���]�����������������������������U��EP�J
����]����������������U��j
j �EP��5����]������������U��EPj
j �MQ�`����]��������U��EP�MQ��A����]������������U��j
j �EP�9����]������������U��EPj
j �MQ�>����]��������U��j
j �EP�25����]������������U��EPj
j �MQ������]��������S�܃������U�k�l$���@�= �}M�C���t�S��K;�t�S���S�݋C��S;�u�C�E���E�    �E��  ��   �Kfn�fE��pE� fE�fpE� fEЋS���  ���  ��   �C�o fE�foE�f�E�fE�foE�fuE�fE�foE�fuE�fE�foE�f�E�fE�foE�f�ȉM��}� t2�U��U��E�C�C�K��C;�u�K�M���E�    �E��:�S���S�*�C��S;�u�C��C���u3���S���S�%�����]��[�������������������������������������������������������������������������������������������������������������SV�L$�T$�\$������tQ+���   t�
:uH��D�B��v4��u�
%�  =�  wً
;u҃�v����������#Ʃ����t�3�^[Íd$ ���^[�����������������������������������������U����=� ��  �} t	�E�   ��E�    �E��E��}� u&hܥh�Yj h�   h��j�
������u̃}� u3��P���    j h�   h��ht�hܥ�%I���������0  �} t	�E�   ��E�    �U�U��}� u&hx�h�Yj h�   h��j�	
������u̃}� u3�JP���    j h�   h��ht�hx��H���������   �}���w	�E�   ��E�    �M�M�}� u&hL�h�Yj h�   h��j�	������u̃}� u0��O���    j h�   h��ht�hL�� H���������.�EP�MQ�UR�������j �EP�MQ�UR�iQ������]�������������������������������������������������������������������������������������������������������������������������U���L�} �n  �EP�M��I���} t	�E�   ��E�    �M��M�}� u#hܥh�Yj j;h��j�D������u̃}� u=�N���    j j;h��h0�hܥ��F�����E�����M��"���E���  �} t	�E�   ��E�    �E��E�}� u#hx�h�Yj j<h��j�������u̃}� u=��M���    j j<h��h0�hx��ZF�����E�����M��!���E��T  �}���w	�E�   ��E�    �U�U�}� u#hL�h�Yj j=h��j�1������u̃}� u=�rM���    j j=h��h0�hL���E�����E�����M�� !���E���   �M���S����   �⃼�    u)�EP�MQ�UR�&�����EЍM�� ���E��   �m�E��M̍M��S��P�U�R�/�����E��E���E�M��UȍM��}S��P�E�P�[/�����E��M���M�U���Ut�}� t�E�;E�t��M�+M��MčM��6 ���E��3���]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�RP�EP�c�����E��}� u	�E�    ��E������E���]�������������������������U���DV�E�    �E�    �E�    jj j �EP�.,�����EĉUȋM�#Mȃ��t#jj j �UR�,�����ẺUЋE�#EЃ��u�
K��� �2  �M+M̋UUЉM܉U��}� �?  
�}� �3  h   j�(P�$�E��}� u%�J���    �E�   �E������E�������   h �  �EP�%�����E�}� |	�}�   r	�E�   ��M܉M��U��U��}� |	�}�   r	�E�   ��E܉E�M�Q�U�R�EP������E��}��u(�	���8u�J���    �E�   �E���EԉU��*�E���M�+ȋE�M܉E��}� �W���|
�}� �K����M�Q�UR��$�����E�Pj �(P��   �}� ��   |
�}� ��   j �MQ�UR�EP�g*�����EԉU؋M�#M؃��t]�UR������P�X��t	�E�    ��E������E虉EԉU؋E�#E؃��u!�*I���    �E�   �� ������0�M�#M؃��t'j �U�R�E�P�MQ��)�����E��U��U�#U����u	��H��� �3�^��]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �}�u�����     �	   �b  �} |�E;<�s	�E�   ��E�    �M��M܃}� u#hhOh�Yj j7h��j�3������u̃}� u;�o���     �iG��� 	   j j7h��h��hhO��?�����	   ��  �E���M������0��D
��t	�E�   ��E�    �M؉Mԃ}� u#hdPh�Yj j8h��j� ������u̃}� u;�����     ��F��� 	   j j8h��h��hdP�&?�����	   �1  �} |�} r	�E�   ��E�    �EЉẼ}� u#h�h�Yj j9h��j� ������u̃}� u;�A���     �;F���    j j9h��h��h��>�����   �   �UR��J�����E�    �E���M������0��D
��t�MQ�UR�EP�5�����E��93�u#h(Nh�Yj jAh��j�Q�������u��E��� 	   �E�	   �E������   ��EP�������ËE�M�d�    Y_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����} t	�E�   ��E�    �E��E��}� u&hp�h�Yj h�   h8�j��������u̃}� u0�HD���    j h�   h8�h��hp��<�����   ��U���3���]���������������������������������������������U����} @  t�} �  t�}   t	�E�    ��E�   �E��E��}� u&h��h�Yj h�   h8�j�2�������u̃}� u0�sC���    j h�   h8�hT�h����;�����   ��U���3���]��������������������������������������������������������U��j�h��h�Ld�    P���SVW���1E�3�P�E�d�    �E�    �} @  t-�} �  t$�}   t�}   t�}   t	�E�    ��E�   �E��E܃}� u#h(�h�Yj j6h8�j��������u̃}� u.�SB���    j j6h8�h��h(��:���������  �}�u�B��� 	   ����  �} |�U;<�s	�E�   ��E�    �E؉Eԃ}� u#hMh�Yj j9h8�j�u�������u̃}� u.�A��� 	   j j9h8�h��hM�:��������2  �U���E������0��T��t	�E�   ��E�    �EЉẼ}� u#h�Mh�Yj j:h8�j���������u̃}� u.�#A��� 	   j j:h8�h��h�M�9��������   �UR��E�����E�    �E���M������0��D
��t�MQ�UR�������E��9�@��� 	   3�u#h(Nh�Yj jEh8�j�4�������u��E������E������   ��UR�������ËE�M�d�    Y_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E���M������0��D
%�   �E��M���U������0��L$�����щU�E�E��}�   $�}�   �a  �}� @  tm�}� �  t$�  �}�   �=  �}�   ��   �  �M���U������0��L������U���E������0��L�`  �E���M������0��D
�   �M���U������0��D�U���E������0��T$�​E���M������0��T$��   �M���U������0��L�ɀ   �U���E������0��L�E���M������0��D
$$��M���U������0��D$�u�U���E������0��T�ʀ   �E���M������0��T�M���U������0��L$�က��U���E������0��L$�}� u� �  ��}� u	� @  ���   ��]�������������������������������������������������������������������������������������������������������������������������������������������������������������U��j�h�d�    P��L���3�P�E�d�    �EP�M�������E�    �} t�M�U��} t	�E�   ��E�    �E��E܃}� u#h��h�Yj j^h��j��������u̃}� uD��;���    j j^h��h<�h���X4�����E�    �E������M�����E��  �} t�}|�}$~	�E�    ��E�   �U؉Uԃ}� u#hP�h�Yj j_h��j��������u̃}� uD�`;���    j j_h��h<�hP��3�����E�    �E������M������E��s  �M�M��E�    �U��E�M���M�M��A����t-�M��A����zt~�M��A��Pj�E�P������E��j�M�Q�M��}A��P�K������EЃ}� t�U��E�M���M���U��-u�E���E�M��U�E���E���M��+u�U��E�M���M�} |�}t�}$~.�} t�U�E��E�    �E������M������E��k  �>�} u8�M��0t	�E
   �&�U����xt�M����Xu	�E   ��E   �} u8�E��0t	�E
   �&�M����xt�E����Xu	�E   ��E   �}u9�U��0u0�E����xt�U����Xu�M���M�U��E�M���M�����3��u�E�j�U�R�M��@��P���������t�E��0�E��Qh  �M�Q�M���?��P��������t0�U��a|�E��z�M�� �M���U�ŰẼ�7�E���f�M�;Mr�\�U���U�E�;E�r�M�;M�u���3��u9U�w�U��UU�U���E���E�} u��M��U�E���E��!����M���M�U��u�} t�E�E��E�    �f�M��u*�U��uV�E��t	�}�   �w�M��u=�}����v4�8��� "   �U��t	�E�������E��t	�E�   ���E�����} t�M�U��E��t�M��ىM�U�U��E������M��o���E��M�d�    Y��]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�EP������]������������������U��j�EP�MQ�UR�EP������]������������������U��=� uj �EP�MQ�URh��L�������j �EP�MQ�URj �0�����]����������������������������U��=� uj�EP�MQ�URh����������j�EP�MQ�URj �������]����������������������������U��EP�MQ�URh�]�
����]�������������������U��EPj �MQh_a������]���������������������U��EP�MQ�URh_a�����]�������������������U��EP�MQ�URhL`�z����]�������������������U��EPj �MQh�]�L����]���������������������U��j�h�h�Ld�    P���SVW���1E�3�P�E�d�    �%���    �� ��E��E�    �} t	�E�   ��E�    �U��U܃}� u#h��h�Yj j4h��j�w�������u̃}� u+�3���    j j4h��h�h���,��������i�M�Q�#�����E�    �U�R������EԋEP�MQ�UR�E�P�U���E؋M�Q�U�R�0�����E������   ��E�P�*����ËE؋M�d�    Y_^[��]���������������������������������������������������������������������������������������U��EPj �MQhL`�����]���������������������U��j�h(d�    P��lVW���3�P�E�d�    �EP�M�������E�    �} t�M�U��} t	�E�   ��E�    �E�E��}� u#h��h�Yj jch@�j��������u̃}� uN��1���    j jch@�h��h���V*�����E�    �E�    �E������M��y���E��U��<  �} t�}|�}$~	�E�    ��E�   �U܉U؃}� u#hP�h�Yj jdh@�j��������u̃}� uN�T1���    j jdh@�h��hP��)�����E�    �E�    �E������M������E��U��  �M�M��E�    �E�    �U��E�M���M�M��7����t-�M��7����zt~�M��7��Pj�E�P�o������E��j�M�Q�M��`7��P�.������Eԃ}� t�U��E�M���M���U��-u�E���E�M��U�E���E���M��+u�U��E�M���M�} u8�U��0t	�E
   �&�E����xt�U����Xu	�E   ��E   �}u9�M��0u0�U����xt�M����Xu�E���E�M��U�E���E�E�RPj�j��P���E��U�j�M�Q�M��[6��P�)�������t�U��0�U��Th  �E�P�M��06��P���������t0�M��a|�U��z�E�� �E���M�MЋUЃ�7�U���   �E�;Er�   �M���M�U�;U�rLw�E�;E�rB�M�;M�u\�U�;U�uT�u�3��E�RPj�j��!���u��}��E��U��E�;E�w,r�M�;M�w"�E�RP�U�R�E�P�b5��3�E�щEȉU���U���U�} u��E��M�U���U�������E���E�M��u�} t�U�U��E�    �E�    �   �E��u:�M��u{�U��t�}�   �w!r�}� w�E��uZ�}����rQw�}��vI�.��� "   �M��t�E������E������&�U��t�E�    �E�   ���E������E�����} t�E�M��U��t�E��؋M̃� �ىEȉM̋UȉU��ẺE��E������M��8���E��U��M�d�    Y_^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��Q�EP�MQ�UR�E�P�������E���]��������������U��=� uj �EP�MQ�URh��,�������j �EP�MQ�URj ������]����������������������������U��j �EP�MQ�UR�EP�������]������������������U��EP�MQ�UR�EP�#����]��������������������U��EP�MQ�UR�9����]��������U��EP�MQ�UR�EP�7#����]��������������������U��=� uj�EP�MQ�URh���������j�EP�MQ�URj � �����]����������������������������U��j�EP�MQ�UR�EP�������]������������������U��EP�MQ�UR�EP�Z�����]��������������������U��EP�MQ�UR�EP�*�����]��������������������U��Q�EPj �MQ�U�R�������E���]����������������U��EP�MQ�UR�P����]��������U��EP�MQ�R����]������������U��EP�MQ�UR�����]��������U��EP�MQ�UR�D����]��������U��EP�MQ�UR�$����]��������U��Q�E�    ��E����E��M���M�U�;Us�E���t�ڋE���]�����������������������U����E�    ���E��M��9 ��   j j j j j��U��Pj j � �E�}� u����   j=h��jj�M�Q�������E��}� u����rj j �U�R�E�Pj��M��Rj j � ��uj�E�P�o���������=j �M�Q���������}�}� tj�U�R�D������E�    �E����E��4���3���]����������������������������������������������������������U��j �EP�MQ�UR� ����]����������������������U���H�EP�M�������} u�E�    �M������E��L  �} t	�E�   ��E�    �M��M��}� u#h8�h�Yj j=h��j��������u̃}� u=��&���    j j=h��h\�h8��O�����E�����M������E���  �} t	�E�   ��E�    �E�E��}� u#h��h�Yj j>h��j�)�������u̃}� u=�j&���    j j>h��h\�h���������E�����M�������E��<  �}���w	�E�   ��E�    �U�U�}� u#h��h�Yj j?h��j��������u̃}� u=��%���    j j?h��h\�h���<�����E�����M��m����E��   �M��a,���H�y u(�UR�EP�MQ�UR�!+�����EЍM��1����E��x�M��(,���@�HQ�UR�EP�MQ�URh  �M��,���@��  Q�M���+��P������ �E�}� u�E�����M�������E���U���UȍM������Eȋ�]������������������������������������������������������������������������������������������������������������������������������������������������������������������U���(�} t�E�M��} t	�E�   ��E�    �U�U�}� u#h��h�Yj j^h��j��������u̃}� u-��#���    j j^h��h�h���J����3��,  �} t�}|�}$~	�E�    ��E�   �M�M��}� u#hP�h�Yj j_h��j�(�������u̃}� u-�i#���    j j_h��h�hP�������3��  �E�E��E�    �M�f�f�U��E����E�j�M�Q�������t�U�f�f�E��M����M����U���-u�E���E�M�f�f�U��E����E���M���+u�U�f�f�E��M����M��} u@�U�R�s ������t	�E
   �&�E����xt�U����Xu	�E   ��E   �}uC�M�Q�- ������u2�U����xt�M����Xu�E����E��M�f�f�U��E����E����3��u�E��M�Q��������E��}��t�V�U���A|	�E���Z~�M���a|9�U���z0�E���a|�M���z�U��� �U���E��E܋M܃�7�M���h�U�;Ur�^�E���E�M�;M�r�U�;U�u���3��u9U�w�E��EE��E���M���M�} u��U�f�f�E��M����M��*����U����U��E��u�} t�M�M��E�    �f�U��u*�E��uV�M��t	�}�   �w�U��u=�}����v4�� ��� "   �E��t	�E�������M��t	�E�   ���E�����} t�U�E���M��t�U��ډU�E��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�UR�:�����]����������������������U��j�EP�MQ�UR�
�����]����������������������U��j �EP�MQ�UR�������]����������������������U��j�EP�MQ�UR������]����������������������U��� �} u#ht�h�Yj jdh�Rj�f�������u̋M�M��U�R�������E��E��H��   u&���� 	   �U��B�� �M��A���  �r  �/�U��B��@t$�Y��� "   �M��Q�� �E��P���  �A  �M��Q��tJ�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J���  ��  �E��H���U��J�E��H���U��J�E��@    �E�    �M�M��U��B%  uC�4���    �� �9E�t� ���    ���9E�u�E�P��������u�M�Q�������U��B%  �  �M��U��+By&h`Sh�Yj h�   h�Rj���������u̋U��E��
+H�M�U��B���M���U��B���M��A�}� ~�U�R�E��HQ�U�R�������E��s�}��t!�}��t�E����M������0��M���E���U��B�� t9jj j �M�Q�V�����E��U�U�#U���u�E��H�� �U��J���  �c�E%��  �M��Qf��*�E�   �E%��  f�E�M�Q�U�R�E�P�d������E��M�;M�t�U��B�� �M��A���  ��E%��  ��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U������3ŉE��N@  f�E�M�    �U�B    �E�@    ��M���M�U���U�} vt�E��M��P�U�@�E��MQ��������UR��������E�P�MQ�������UR�������E��M��E�    �E�    �U�R�EP�������t����M�y uB�U�B���M�A�U�B���M���M�A�U����M��U��f�U�뵋E�H�� �  u�UR�-�����f�E�f��f�E��؋Mf�U�f�Q
�M�3��]�����]�������������������������������������������������������������������������������������������������U��j�hXd�    P��pVW���3�P�E�d�    �EP�M�������E�    �} t�M�U��} t	�E�   ��E�    �E�E��}� u#h��h�Yj jch�j��������u̃}� uN�����    j jch�h|�h���F�����E�    �E�    �E������M��i����E��U��P  �} t�}|�}$~	�E�    ��E�   �U܉U؃}� u#hP�h�Yj jdh�j��������u̃}� uN�D���    j jdh�h|�hP�������E�    �E�    �E������M�������E��U��  �M�M��E�    �E�    �U�f�f�E��M���M�j�U�R��������t�E�f�f�M��U���U����E���-u�M���M�U�f�f�E��M���M���U���+u�E�f�f�M��U���U�} |�}t�}$~8�} t�E�M��E�    �E�    �E������M�������E��U���  �F�} u@�U�R���������t	�E
   �&�E����xt�U����Xu	�E   ��E   �}uC�M�Q��������u2�U����xt�M����Xu�E���E�M�f�f�U��E���E�E�RPj�j��#����EĉU��M�Q�>������E�}��t�Y�U���A|	�E���Z~�M���a|9�U���z0�E���a|�M���z�U��� �U���E��EԋMԃ�7�M���   �U�;Ur�   �E���E�M�;M�rLw�U�;U�rB�E�;E�u\�M�;M�uT�u�3��E�RPj�j�������u��}��E��U��U�;U�w,r�E�;E�w"�E�RP�M�Q�U�R�@��3�E�щẺU���U���U�} u��E�f�f�M��U���U�������E���E�M��u�} t�U�U��E�    �E�    �   �E��u:�M��u{�U��t�}�   �w!r�}� w�E��uZ�}����rQw�}��vI����� "   �M��t�E������E������&�U��t�E�    �E�   ���E������E�����} t�E�M��U��t�E��؋MЃ� �ىẺMЋỦU��EЉE��E������M������E��U��M�d�    Y_^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    j j j j j��EPj j � �E��}� u�� P�&���������   h�  h��j�M�Q�U������E��}� u���   j j �U�R�E�Pj��MQj j � ��u!�� P�������j�U�R���������X�E�    �E�P�MQ�U�R�E�P��������} t"�}� t�M�+M��U�J�M��	�U�    j�E�P�.������E���]������������������������������������������������������������������������U��=� uj �EP�MQ�URh����������j �EP�MQ�URj �������]����������������������������U��j �EP�MQ�UR�EP������]������������������U��EP�MQ�UR�EP�������]��������������������U��EP�MQ�UR�1�����]��������U��EP�MQ�UR�EP������]��������������������U��=� uj�EP�MQ�URh����������j�EP�MQ�URj �������]����������������������������U��j�EP�MQ�UR�EP������]������������������U��EP�MQ�UR�EP�������]��������������������U��EP�MQ�UR�EP������]��������������������U��j �EP�MQ������]����������U��EP�MQ�UR������]��������U��EP�MQ�a�����]������������U��EP�MQ�UR�n�����]��������U��EP�MQ�UR������]��������U��EP�MQ�UR������]��������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_���������������������������������U���\���3ŉE��E�E��MQ�M������} t�U�E��} t	�E�   ��E�    �MȉMă}� u#h��h�Yj jDh��j��������u̃}� u;�����    j jDh��h,�h���.�������]��M��a����E��B  �M��U����t/�M��I��� �xt~�M��9��Pj�M��R�"������E��j�E��Q�M����P��������Eԃ}� t�U����U�뗍M�����P�E�P�M�Q�������E܃} t�U܋E�B�M��U܋�E؋M؁�@  t���]̃} t�U�E��p�M؁�   t.�U����-u������]��	����]����� "   �7�M؁�   t#�U��B��������Dz���]��{��� "   �	�E��@�]��E��]��M������E��M�3��������]�������������������������������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�������]����������U���0V�E�    �E�    �} t	�E�   ��E�    �E܉E؃}� u#hD�h�Yj jShp�j���������u̃}� u.�<���    j jShp�h��hD����������  �U��E�}� tj=�M�Q�������E��}� t�U�;U�u��
���    ����A  �E�+E�=�  |#h��h�Yj jehp�j�W�������u�h�  �U���R�����=�  r#h0�h�Yj jfhp�j��������u̋M��Q��u	�E�   ��E�    �EԉE� �;��u� �R��  ��� ��= � ��   �} t*�=� t!�w����t��	���    ����X  �   �}� t3��F  �   �= � u7h�   h��jj脿����� ��= � u����  � ��     �=� u8h�   h��jj�D��������=� u�����  ���    � ��U��}� u23�u&h��h�Yj h�   hp�j���������u̃���  �U�+U�R�E�P�0  ���E��}� ��   �M��9 ��   j�U��E���Q� ������}� ti�	�U����U��E��M��<� t�U��E��M��u��L����ց}����?s2h�   h��jj�U�R� �P��	�����E��}� t	�M�� ���U��E��M���U�    �   �}� ��   �}� }�E��؉E��M���;M�|;�U��������?s-h�   h��j�E���Pj� �Q�^	�����E��}� u����P  �U��E��M���U��E��D�    �M�    �U�� ��j�E�P��������M�    3��  �} ��   h  h��jj�U�R�P�������P�������E�}� ��   j h  hp�h��h ��E�P�M�Q��������P�U�R�\����P�������E�+E�E�E�M�� �U���U�}� t	�E�    ��E�EЋM�Q�U�R�\��u�E������}��u����� *   j�E�P�������}� tj�M�Q��������U�    �E�^��]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����E�    �E�E��} u3���   �M���U�E����E��}� t�M���M���h�  h��jj�U��R�������E��E��E�}� u
j	�0������M�M��U��: ��   �E��Q���������E�h�  h��jj�U�R�������M���U��: t7j h�  hp�h��h���E��Q�U�R�E��Q�����P��������U����U��E����E��k����M��    �E��]������������������������������������������������������������������������������U��Q� ��E��	�M����M��U��: tK�EP�M��R�EP���������u/�M���E���=t�U���M���u�E�+ ����뤋E�+ ����؋�]�������������������������������������U��=� u�EP�MQ�UR�>�������j �EP�MQ�UR�����]���������������������U���H�EP�M��C����} u�E�    �M��x����E��q  �} t	�E�   ��E�    �M��M��}� u#h h�Yj j?h@ j�!�������u̃}� u=�b���    j j?h@ h� h �������E�����M�������E���  �} t	�E�   ��E�    �E�E��}� u#h� h�Yj j@h@ j虻������u̃}� u=�����    j j@h@ h� h� �7������E�����M��h����E��a  �}���w	�E�   ��E�    �U�U�}� u#hL�h�Yj jAh@ j��������u̃}� u=�O���    j jAh@ h� hL��������E�����M�������E���   �M�������   �� ���    u0�M����P�EP�MQ�UR�������EЍM������E��   �M����� �HQ�UR�EP�MQ�URh  �M��b��� �   �� ���   R�M��H��P�N����� �E�}� u�o ���    �E�����M������E���E���EȍM������Eȋ�]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���E��0}����
  �M��:}�E��0��  �U���  ��  �E=`  }�����  �M��j  }�E-`  �  �U���  }����  �E=�  }�E-�  �  �M��f	  }����w  �U��p	  }�E-f	  �]  �E=�	  }����J  �M���	  }�E-�	  �0  �U��f
  }����  �E=p
  }�E-f
  �  �M���
  }�����  �U���
  }�E-�
  ��  �E=f  }�����  �M��p  }�E-f  �  �U��f  }����  �E=p  }�E-f  �{  �M���  }����g  �U���  }�E-�  �M  �E=f  }����:  �M��p  }�E-f  �   �U��P  }����  �E=Z  }�E-P  ��   �M���  }�����   �U���  }�E-�  ��   �E=   }����   �M��*  }�E-   �   �U��@  }����   �E=J  }�E-@  �n�M���  }����]�U���  }�E-�  �F�E=  }����6�M��  }�E-  ������U���  }�E-�  ����]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���X���3ŉE��E�E��MQ�M������} t�U�E��} t	�E�   ��E�    �MЉMԃ}� u#h��h�Yj jGh� j��������u̃}� u;�!����    j jGh� hTh���~��������]��M������E���   j�E��Q���������t�U����U����M����P�E�P�M�Q��������E܃} t�U܋B�M��A�E��M܋�U؋E�%@  t���]ȃ} t�M�U��n�E�%�   t.�M����-u������]��	����]��A���� "   �6�E�%   t#�M��A��������Dz���]������ "   �	�U��B�]��E��]��M������E��M�3��`�����]��������������������������������������������������������������������������������������������������������������������U��j �EP�MQ�������]����������U���(���3ŉE��E�    �EPj j j j �MQ�U�R�E�P������ �E�M��t�U��   �U��E�    �E�    �F�E�P�M�Q�:������E�U��u�}�u�E��   �E�M��u�}�u�U��   �U�E�M��U�+U�E�P�M�U܉Q�E��A�E�M�3��������]���������������������������������������������������������U��j �EP�MQ�U�����]����������U���4�EP�M�胻���} t	�E�   ��E�    �M��M�}� u#hlh�Yj j:h�j�~�������u̃}� u=�����    j j:h�h�hl�������E�    �M��M����E���   �M��A����@�x u#�MQ�UR��������E�M������E���   �	�E���E�Mf�f�U��E���t|�M�������H�U��D��tS�M���M�U���u�E�    �M������E��j�M����U��9Mu�M���M�M������E��@��U�9Uu��h����E�9Eu�M�M��M��`����E���E�    �M��L����E܋�]�������������������������������������������������������������������������������������������������������U���(���3ŉE��E�    �EPj j j j �MQ�U�R�E�P�%����� �E�M��t�U��   �U��E�    �E�    �F�E�P�M�Q�
������E�U��u�}�u�E��   �E�M��u�}�u�U��   �U�E�M��U�+U���E�P�M�U܉Q�E��A�E�M�3��������]������������������������������������������������������̃= �r_�D$�����fn��p� ۋT$�   ���#���+��o
f��ft�ft�f��f��#�u����������f~�3�:E��3��D$S�����T$��   t�
��:�tY��tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u!% �t�% u��   �u�^_[3�ÍB�[ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��������������������������������������������������������������������������������������U������3ŉE��EPj j j �MQ�UR�EP�M�Q������ �E�UR�E�P�/������E�}�u	�M���M�E�M�3�������]�����������������������������������������U���   ���3ŉE��E��E�3�f�M�ǅl���   �E�    �E�    �E�    ǅp���    �E�    ǅ|���    �E�    �E�    �E�    �E�    3�f�U�3�f�E��E�    �E�    �}$ tǅh���   �
ǅh���    ��h�����\�����\��� u#h��h�Yj j~h�j�ҫ������u̃�\��� u-�����    j j~h�hh���m�����3���  �E�E̋M̉M��	�Ũ��ŰE���� t!�U����	t�M����
t�E����u�Ƀ}�
�N  �U�f�f�EЋM̃��M̋Uȉ�`�����`����   ��`����$�̂�MЃ�1|�UЃ�9�E�   �Ẽ��E��   �MЋU$����   ��;�u	�E�   �a�EЉ�t�����t���+t��t���-t#��t���0t�*�E�   �1�E�   3�f�M��"�E�   � �  f�U���E�
   �Ẽ��E��e  �E�   �MЃ�1|�UЃ�9�E�   �Ẽ��E��|�MЋU$����   ��;�u	�E�   �[�EЉE��M���+�M��}�:w5�U�����$����E�   �+�E�   �"�M̃��M��E�   ��E�
   �Ũ��U��  �EЃ�1|�MЃ�9�E�   �Ũ��U��L�EЋM$����   ��
;�u	�E�   �+�UЉ�T�����T���0t�	�E�   ��E�
   �E��E��D  �E�   ��M�f�f�UЋẼ��E��MЃ�0|:�UЃ�91�}�s �E����E��MЃ�0�U��
�E����E��	�M����M���UЋE$����   ��;�u	�E�   �R�MЉM��U���+�U��}�:w,�E���T��$�H��E�   �"�Ũ��U��E�   ��E�
   �Ẽ��E��m  �E�   �E�   �}� u)��M�f�f�UЋẼ��E��MЃ�0u�U����U�����E�f�f�MЋŨ��U��EЃ�0|8�MЃ�9/�}�s'�U����U��EЃ�0�M���U����U��E����E���MЉM��U���+�U��}�:w,�E������$����E�   �"�Ũ��U��E�   ��E�
   �Ẽ��E��  �E�   �MЃ�0|�UЃ�9�E�   �Ẽ��E���E�
   �M��M��F  �Ũ��U��EЃ�1|�MЃ�9�E�	   �Ũ��U��Y�EЉ�x�����x���+t0��x���-t��x���0t�%�E�   �)�E�   ǅl���������E�   ��E�
   �M��M��  ǅp���   ��U�f�f�EЋM̃��M��UЃ�0u���EЃ�1|�MЃ�9�E�	   �Ũ��U���E�
   �Ẽ��E��X  �MЃ�1|�UЃ�9�E�	   �Ẽ��E��+�MЉ�X�����X���0t�	�E�   ��E�
   �U��U��  ǅp���   �E�    ��E�f�f�MЋŨ��U��EЃ�0|,�MЃ�9#kU�
�EЍLЉM��}�P  ~	�E�Q  �븋U��U���E�f�f�MЋŨ��U��EЃ�0|�MЃ�9���E�
   �Ũ��U��h�}  tR�Ẽ��E��MЉ�d�����d���+t��d���-t��E�   ǅl���������E�   ��E�
   �U��U���E�
   �Ẽ��E������M�Ủ�}� �`  �}� �V  ��|��� �I  �}�vF�   k��T���|�   k��T����   k��T��E�   �U����U��E����E��}� ��   �M����M��	�U����U��E����u�U����U��E����E��ٍM�Q�U�R�E�P�A�������l��� }�M��ىM��U�U��U���p��� u	�E�E�E��}� u	�M�+M�M��}�P  ~	�E�   �E�}�����}ǅ|���   �0�UR�E�P�M�Q�.�����f�U�f�U��E։E��MډM�f�U�f�U��3�f�E�3�f�M��UĉU��E��E��}� u$3�f�M�3�f�U��EĉE��M��M��U����U��Y�}� t(��  f�E��E�   ��E�    3�f�M��U����U��+��|��� t"3�f�E�3�f�M��UĉU��E��E��M����M��Uf�E�f��M�U��Q�E�M��H�U��E�ЋMf�Q
�E��M�3�������]ÍI ~z,{�{M|$}~K~9�~���)��{�{�{�{  ��|�|}  ��}�}�}  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%  �% �% �% �% �% �% �% �%  �%$ �%( �%, �%0 �%4 �%8 �%< �%@ �%D �%H �%L �%P �%T �%X �%\ �%` �%d �%h �%l �%p �%t �%x �%| �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �%� �% �%�%�%�%�%�%�%�% �%$�%(�%,�%0�%4�%8�%<�%@�%D�%H�%L�%P�%T�%X�%\�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋T$�B�� ���3�������;���������������������̋T$�B�� ���3������(<�ܦ�������������������̋T$�B������3�资���;鬦�������������������̋T$�B������3�腄���J�3��{����X9�r��������������������������̋T$�B������3��E����J�3��;�����9�2��������������������������̋T$�B�� ���3�������:����������������������̋T$�B������3��Ճ���h;�̥�������������������̋T$�B������3�襃���J�3�蛃���H:钥�������������������������̋M��2w���M���� ����T$�B�J�3��U�����@�L��������������������̋M���v���T$�B�J�3�� ����d@�����������������j8h�o�E�P�E�P�(s����ËT$�B�J�3��������?�פ��������������̍M�锛��h���E�P��m����ËT$�B�J�3�螂����@镤����������������������������̍M��D����T$�B�J�3��`����4@�W����������������h�   h�o�E�P�E�P�Rl����ËT$�B�J�3������@������������������������������h�   h�o�E�P�E�P�l����ËT$�B�J�3��́����?�ģ���������������������������̍M���p���T$�B�J�3�萁���J�3�膁����G�}���������������������̍M��4����T$�B�J�3��P�����D�G���������������̍M������T$�B�J�3�� ����lF����������������̍M��ԙ���T$�B�J�3�������pG����������������̋M��t���T$�B�J�3�������LB鷢��������������̋M��bt���T$�B�J�3�萀���hE釢��������������̋M��2t���T$�B�J�3��`�����F�W���������������̍�`�����]���M��jo����p�����]���M��Wo���T$�B��0���3������J�3�������E���������������������������������������h  h���E�P�E�P��i����ËE����   �e���M��]���ËT$�B�J�3�����B鋡�����������������������������������hD  h���E�P�E�P�ri����ËE����   �e���M�����ËT$�B�J�3��$���4E�������������������������������������h�   h���E�P�E�P�i����ËE����   �e���M��}���ËT$�B�J�3��~����F髠����������������������������������̍�\����7\���M��m����`����$\���M��m���T$�B��`���3��O~���J�3��E~���tD�<������������������������������������̍�P�����[���M��:m����T����[���M��'m���T$�B��T���3���}���J�3���}����D�̟�����������������������������������̍M���l���M���l���T$�B��X���3��}���J�3��{}���(D�r��������������������������̋T$�B��l���3��E}���J�3��;}���<G�2��������������������������̍M���Z���M��=l���M��Z���M��-l���T$�B��L���3���|���J�3���|���8F�Ҟ�������������������������̍M�鄕���T$�B�J�3��|���A闞��������������̍M��8����M��L����T$�B�J�3��h|���DA�_������������������������jJhȂ�E�P�E�P�Uf�����jKhȂ�E�P�E�P�=f�����jLhȂ�E�P�E�P�%f�����jMhȂ�E�P�E�P�f�����jOhȂ�E�P�E�P��e����ËT$�B�J�3���{���pA鷝����������������������������������������������̍M��:Y���T$�B�J�3��p{���J�3��f{����B�]���������������������̍M���X���T$�B�J�3��0{���J�3��&{��� C����������������������̍M��X���T$�B�J�3���z���J�3���z���0C�ݜ��������������������̍M��zX���T$�B�J�3��z���J�3��z���`C靜��������������������̍M��:X���T$�B�J�3��pz���J�3��fz����C�]���������������������̍M���W���T$�B�J�3��0z���J�3��&z����C����������������������̍M��W���T$�B�J�3���y���J�3���y����C�ݛ��������������������̍�H����wW���M���h����|�����h���M���h����`����QW���T$�B��@���3��y���J�3��zy���tB�q�������������������������̍�p����W���M��zh���T$�B��d���3��2y���J�3��(y����E������������������������̍M��V���M��̑���T$�B�J�3���x����A�ߚ����������������������̍M���g���T$�B�J�3��x���J�3��x����q靚��������������������̍M��g���T$�B�J�3��px���J�3��fx����p�]���������������������̍M��ug���T$�B�J�3��0x���J�3��&x���(q����������������������̍M��5g���T$�B�J�3���w���J�3���w����p�ݙ��������������������̍M��]���M�]���M��]���M��]���M��]���M���]���M��]���T$�B�J�3��w����r�w�������������������������������̍M�e���M�e���M��e���M��e���M��e���M���R���M��e���T$�B�J�3��w���r��������������������������������̋EP�E�P�(b����ËT$�B�J�3���v���8s龘���������������������̋EP�E�P��a����ËT$�B�J�3��v���s�~����������������������̍M��4����T$�B�J�3��Pv����o�G���������������̍M������T$�B�J�3�� v���p]����������������̍M��Ԏ���T$�B�J�3���u��� d����������������̍M�餎���T$�B�J�3���u���,U鷗��������������̍M��t����T$�B�J�3��u���8K釗��������������̍M��D����T$�B�J�3��`u���K�W���������������̍M������T$�B�J�3��0u����d�'���������������̍M������T$�B�J�3�� u����U�����������������̍M�鴍���T$�B�J�3���t����f�ǖ��������������̍M�鄍���T$�B�J�3��t����W闖��������������̍M��T����T$�B�J�3��pt����j�g���������������̍M��$����T$�B�J�3��@t����Y�7���������������̍M������T$�B�J�3��t���hl����������������̍M��Č���T$�B�J�3���s����k�ו��������������̍M�锌���T$�B�J�3��s���[駕��������������̍M��d����T$�B�J�3��s����Z�w���������������̍M��4����T$�B�J�3��Ps����`�G���������������̍M������T$�B�J�3�� s����Q����������������̍M��ԋ���T$�B�J�3���r���b����������������̍M�餋���T$�B�J�3���r���0S鷔��������������̍M��t����T$�B�J�3��r���c釔��������������̍M��D����T$�B�J�3��`r���4T�W���������������̍M������T$�B�J�3��0r���\n�'���������������̍M������T$�B�J�3�� r���]�����������������̍M�鴊���T$�B�J�3���q���xo�Ǔ��������������̍M�鄊���T$�B�J�3��q���@]闓��������������̋M��jV���T$�B�J�3��pq��� k�g���������������̋M��:V���T$�B�J�3��@q����Y�7���������������̋M��Y���T$�B�J�3��q���Hh����������������̋M���P���T$�B�J�3���p���hK�ג��������������̋M�������T$�B�J�3��p����p駒��������������̋M�鏁���T$�B�J�3��p����o�w���������������̋M��_T���T$�B�J�3��Pp���xh�G���������������̋M��/T���T$�B�J�3�� p���8i����������������̋M���S���T$�B�J�3���o���i����������������̋M���S���T$�B�J�3���o����h鷑��������������̋M��S���T$�B�J�3��o����h金��������������̋M��#Y���T$�B�J�3��`o����K�W���������������̋M���X���T$�B�J�3��0o���XL�'���������������̋M���X���T$�B�J�3�� o���(L�����������������̋M��X���T$�B�J�3���n����K�ǐ��������������̋M��cX���T$�B�J�3��n����K闐��������������̋M���p���T$�B�J�3��pn����I�g���������������̋M��p���T$�B�J�3��@n���8I�7���������������̋M���a���T$�B�J�3��n���8c����������������̋M��a���T$�B�J�3���m���dT�׏��������������̋M���U���T$�B�J�3��m����J駏��������������̋M��U���T$�B�J�3��m��� J�w���������������̋M��{���T$�B�J�3��Pm���0d�G���������������̋M��{���T$�B�J�3�� m���\U����������������̋M���`���T$�B�J�3���l����d����������������̋M��`���T$�B�J�3���l��� V鷎��������������̋M��b`���T$�B�J�3��l����f野��������������̋M��2`���T$�B�J�3��`l����W�W���������������̋M��`���T$�B�J�3��0l����]�'���������������̋M���_���T$�B�J�3�� l���O�����������������̋M��_���T$�B�J�3���k��� a�Ǎ��������������̋M��r_���T$�B�J�3��k���,R闍��������������̋M��B_���T$�B�J�3��pk���4b�g���������������̋M��_���T$�B�J�3��@k���`S�7���������������̋M��Đ���T$�B�J�3��k����l����������������̋M�锐���T$�B�J�3���j���L[�׌��������������̋M��^���M����$����T$�B�J�3��j����n霌�������������������̋M��B^���M��������T$�B�J�3��ej����M�\��������������������̍M��GP���T$�B�J�3��0j����q�'���������������̍M��bP���T$�B�J�3�� j����q�����������������̍M��HX���T$�B�J�3���i���8p�ǋ��������������̍M��E���T$�B�J�3��i���hp闋��������������̍M��O���T$�B�J�3��pi���Xq�g���������������̍M��W���T$�B�J�3��@i���p�7���������������̋T$�B�J�3��i��� j������������������������̋T$�B�J�3���h���@M�ߊ����������������������̍�`����wF���M��Y����p����dF���M���W���T$�B��0���3��h���J�3��h����a�|������������������������������������̍�`����F���M��u����p�����E���M��gW���T$�B��0���3��h���J�3��h����R��������������������������������������h^  h��E�P�E�P��Q����ËE����   �e���M��m���ËT$�B�J�3��g����I雉�����������������������������������hs  h��E�P�E�P�Q����ËE����   �e���M������ËT$�B�J�3��4g���xI�+������������������������������������jChX��E�P�E�P�Q����ËEЃ��   �e���M��V��ËEЃ��   �e����|����t���ËT$�B�J�3��f���J�3��f���`c阈��������������������������������jChX��E�P�E�P�P����ËEЃ��   �e���M��}U��ËEЃ��   �e����|�������ËT$�B�J�3��f���J�3��f����T����������������������������������hO  h��E�P�E�P��O����ËE����   �e���M��m���ËT$�B�J�3��e����J雇�����������������������������������hl
  h��E�P�E�P�O����ËE����   �e���M������ËT$�B�J�3��4e���`J�+������������������������������������jMh��E�P�E�P�O����ËE����   �e���M�鐏��ËT$�B�J�3���d���pd龆����������������������jMh��E�P�E�P�N����ËE����   �e���M��0���ËT$�B�J�3��gd����U�^�����������������������h�  h��E�P�E�P�RN����ËE����   �e���M��͎��ËT$�B�J�3��d���e��������������������������������������h�  h��E�P�E�P��M����ËE����   �e���M��]���ËT$�B�J�3��c���@V鋅�����������������������������������h�  h��E�P�E�P�rM����ËE����   �e���M�����ËT$�B�J�3��$c����f�������������������������������������h�  h��E�P�E�P�M����ËE����   �e���M��}���ËT$�B�J�3��b���X髄�����������������������������������h(  h��E�P�E�P�L����ËE����   �e���M�����ËT$�B�J�3��Db���4l�;������������������������������������h(  h��E�P�E�P�"L����ËE����   �e���M�靌��ËT$�B�J�3���a����k�˃�����������������������������������h(  h��E�P�E�P�K����ËE����   �e���M��-���ËT$�B�J�3��da����Z�[������������������������������������h(  h��E�P�E�P�BK����ËE����   �e���M�齋��ËT$�B�J�3���`���tZ�������������������������������������h  h���E�P�E�P��J����ËE����   �e���M��M���ËT$�B�J�3��`����]�{������������������������������������h  h���E�P�E�P�bJ����ËE����   �e���M��݊��ËT$�B�J�3��`����N�������������������������������������hD  h���E�P�E�P��I����ËE����   �e���M��m���ËT$�B�J�3��_����`雁�����������������������������������hD  h���E�P�E�P�I����ËE����   �e���M������ËT$�B�J�3��4_����Q�+������������������������������������h�   h���E�P�E�P�I����ËE����   �e���M�鍉��ËT$�B�J�3���^���tb黀�����������������������������������h�   h���E�P�E�P�H����ËE����   �e���M�����ËT$�B�J�3��T^����S�K������������������������������������h�   h���E�P�E�P�2H����ËE����   �e���M�魈��ËT$�B�J�3���]����l�������������������������������������h�   h���E�P�E�P��G����ËE����   �e���M��=���ËT$�B�J�3��t]����[�k�����������������������������������h  h���E�P�E�P�RG����ËE����   �e���M��͇��ËT$�B�J�3��]����n��~�����������������������������������h|  h���E�P�E�P��F����ËE����   �e���M��]���ËT$�B�J�3��\���,N�~����������������������������������̍�L����:���M��K����P����:���M��wK���T$�B��P���3��/\���J�3��%\���`�~�����������������������������������̍�L����9���M��K����P����9���M��K���T$�B��P���3��[���J�3��[���8Q�}�����������������������������������̍�0����79���M��J����4����$9���M��J���T$�B��4���3��O[���J�3��E[���X`�<}�����������������������������������̍�0�����8���M��:J����4����8���M��'J���T$�B��4���3���Z���J�3���Z����Q��|�����������������������������������̍M��Z8���T$�B�J�3��Z���,n�|��������������̍M��*8���T$�B�J�3��`Z����\�W|��������������̍M��uI���M��mI���T$�B��8���3��%Z���J�3��Z����_�|�������������������������̍M��%I���M��I���T$�B��8���3���Y���J�3���Y����P��{�������������������������̍������W7���������L7���M���I���M��H���������17���M��I��������?����h����`?����|������   ��|������\����??��Í�D����3?����|������   ��|�����������XI��Ë�|������   ��|�����������6I��Ë�|������   ��|����������I��Ë�|������   ��|���������H��Í�d�����G���M���G����������>����,����>����|����� �   ��|���ߍ�P����a>��Í�8����U>���T$�B��0���3��;X���J�3��1X����e�(z���������������������������������������������������������������������������������������������������������������̍������g5���������\5���M��fd���M���F���������A5���M��Kd��������D3����h�����E����|������   ��|������\����E��Í�D����E����|������   ��|������������c��Ë�|������   ��|������������c��Ë�|������   ��|����������c��Ë�|������   ��|��������c��Í�d�����E���M���E���������f2����,�����D����|����� �   ��|���ߍ�P�����D��Í�8�����D���T$�B��0���3��KV���J�3��AV����V�8x���������������������������������������������������������������������������������������������������������������̋T$�B�J�3��U���J�3��U���|k�w������������̋T$�B�J�3��U���J�3��~U���0Z�uw������������̋T$�B��l���3��UU���J�3��KU����b�Bw�������������������������̋T$�B��l���3��U���J�3��U��� T�w�������������������������̋T$�B�J�3���T���8m��v����������������������̋T$�B�J�3��T����[�v����������������������̍M���|���T$�B�J�3��pT���o�gv��������������̍M��|���T$�B�J�3��@T���`N�7v��������������̍M���1���M��eD���M���1���M��=C���T$�B��L���3���S���J�3���S����a��u�������������������������̍M��z1���M��`���M��j1���M���B���T$�B��L���3��S���J�3��S����R�u��������������������������jUh��E�P�E�P�u=�����jVh���P���P�E�P�Z=�����jWh���8���P�E�P�?=�����jXh���H���P�E�P�$=�����jYh���(���P�E�P�	=�����jZh���@���P�E�P��<�����j[h���0���P�E�P��<�����j\h���|���P�E�P�<�����j]h���l���P�E�P�<�����j^h���\���P�E�P�<�����j_h���L���P�E�P�g<�����j`h���<���P�E�P�L<�����jbh���,���P�E�P�1<����ËT$�B��,���3���Q���dH��s��������������������������������������������������������������������������������������������������������j-h��E�P�E�P�;�����j.h���P���P�E�P�z;�����j/h���8���P�E�P�_;�����j0h���H���P�E�P�D;�����j1h���(���P�E�P�);�����j2h���@���P�E�P�;�����j3h���0���P�E�P��:�����j4h���|���P�E�P��:�����j5h���l���P�E�P�:�����j6h���\���P�E�P�:�����j7h���L���P�E�P�:�����j8h���<���P�E�P�l:�����j:h���,���P�E�P�Q:����ËT$�B��,���3��P����G�r�������������������������������������������������������������������������������������������������������̍M��5���M��5���T$�B�J�3��O����j�q����������������������̍M�0+���M�(+���T$�B�J�3��HO����M�?q����������������������̍M�r5���T$�B�J�3��O����j�q��������������̍M��*���T$�B�J�3���N���tY��p��������������̍M$�?���������o,����t����d,���M���=���M���>���M���>��������4����$����4��������x4���������m4���������b4���������W4���������L4���������A4���� ����64���T$�B��t���3��N���J�3��N����g�	p����������������������������������������������������������������̍M$�Z���������o+����t����d+���M���<���M��fZ���M��^Z���������;����$�����;���������;����������;����������;���������;���������;���������;���� ����;���T$�B��t���3��M���J�3��M����X�	o����������������������������������������������������������������̍M���;���T$�B�J�3��L���J�3��L���He�n��������������������̍M��;���T$�B�J�3��pL���J�3��fL���xe�]n��������������������̍M��u;���T$�B�J�3��0L���J�3��&L���tV�n��������������������̍M��5;���T$�B�J�3���K���J�3���K����V��m��������������������̍M��z)���T$�B�J�3��K���J�3��K���h^�m��������������������̍M��:)���T$�B�J�3��pK���J�3��fK����^�]m��������������������̍M���(���T$�B�J�3��0K���J�3��&K����^�m��������������������̍M��(���T$�B�J�3���J���J�3���J����^��l��������������������̍M��z(���T$�B�J�3��J���J�3��J����_�l��������������������̍M��:(���T$�B�J�3��pJ���J�3��fJ���(_�]l��������������������̍M���'���T$�B�J�3��0J���J�3��&J���X_�l��������������������̍�H����'���M��B:����|����7:���M��/:����`����'���T$�B��@���3���I���J�3��I���^�k������������������������̍M��J'���T$�B�J�3��I���J�3��vI����O�mk��������������������̍M��
'���T$�B�J�3��@I���J�3��6I����O�-k��������������������̍M���&���T$�B�J�3�� I���J�3���H����O��j��������������������̍M��&���T$�B�J�3���H���J�3��H���$P�j��������������������̍M��J&���T$�B�J�3��H���J�3��vH����P�mj��������������������̍M��
&���T$�B�J�3��@H���J�3��6H���TP�-j��������������������̍M���%���T$�B�J�3�� H���J�3���G����P��i��������������������̍�H����%���M��T����|����T���M��~T����`����a%���T$�B��@���3��G���J�3��G���8O�i������������������������̍M��%���T$�B�J�3��PG����m�Gi��������������̍M���$���T$�B�J�3�� G����\�i��������������̍M��$���T$�B�J�3���F����m��h��������������̍M��$���T$�B�J�3���F���P\�h��������������̍M��Z$���T$�B�J�3��F���lm�h��������������̍M��*$���T$�B�J�3��`F��� \�Wh��������������̍M���#���T$�B�J�3��0F����m�'h��������������̍M���#���T$�B�J�3�� F����\��g��������������̍M��#���M��%6���T$�B�J�3���E���J�3��E���hg�g����������������������������̍M��J#���M���5���T$�B�J�3��xE���J�3��nE���,g�eg����������������������������̍M���"���M��R���T$�B�J�3��(E���J�3��E����X�g����������������������������̍M��"���M��Q���T$�B�J�3���D���J�3���D���XX��f����������������������������̍�p����W"���M���4���T$�B��d���3��D���J�3��xD���8a�of����������������������̍�p����"���M��Q���T$�B��d���3��2D���J�3��(D���dR�f����������������������̍M���P���M��`2���T$�B�J�3���C���J�3���C���Do��e����������������������������̍M��|P���M��2���T$�B�J�3��C���J�3��C����N�e����������������������������̍M��3���M��_)���M��W)���T$�B�J�3��@C���J�3��6C����c�-e��������������������̍M���O���M��p1���M��h1���T$�B�J�3���B���J�3���B����T��d��������������������̋E����   �e���M���1��ËT$�B�J�3��B���J�3��B���I�d�������������������̍M,�w(���M �o(���M�(���M�(���M��(����p����L(���M��(����|����(����d����.(���M��q(���T$�B��l���3��B���`i�d������������������������������������������̍M,�80���M �00���M����M����M������p����0���M��m����|����b����d�����/���M��O���T$�B��l���3��lA����L�cc������������������������������������������̍M�C>���M�;>���M��3>���M��+>���M��#>���M��,(���M��>���T$�B�J�3���@���D��b������������������������������̍M��Y���T$�B�J�3��@����u�b��������������̍M��dY���T$�B�J�3��@���0v�wb��������������̍M��4Y���T$�B�J�3��P@���x�Gb��������������̍M��Y���T$�B�J�3�� @���z�b��������������̍M���X���T$�B�J�3���?���|{��a��������������̍M��X���T$�B�J�3���?���{�a��������������̍M��tX���T$�B�J�3��?���p}�a��������������̍M��DX���T$�B�J�3��`?����~�Wa��������������̋M��*$���T$�B�J�3��0?���4z�'a��������������̋M���D���T$�B�J�3�� ?���hs��`��������������̋M��2���T$�B�J�3���>����t��`��������������̋M��M���T$�B�J�3��>����u�`��������������̋M��B2���T$�B�J�3��p>���`v�g`��������������̋M��2���T$�B�J�3��@>���<x�7`��������������̋M���c���T$�B�J�3��>����{�`��������������̋M��1���M����Tf���T$�B�J�3���=����}��_�������������������̍M���:���T$�B�J�3��=����~�_��������������̍M��$���T$�B�J�3��p=����g_��������������̍M��c:���T$�B�J�3��@=����~�7_���������������jChX��E�P�E�P�5'����ËEЃ��   �e���M��-,��ËEЃ��   �e����|����g��ËT$�B�J�3���<���J�3���<����t�^��������������������������������jMh��E�P�E�P�&����ËE����   �e���M�� g��ËT$�B�J�3��W<����u�N^����������������������h�  h��E�P�E�P�B&����ËE����   �e���M��f��ËT$�B�J�3���;����v��]�����������������������������������h�  h��E�P�E�P��%����ËE����   �e���M��Mf��ËT$�B�J�3��;���|x�{]�����������������������������������h(  h��E�P�E�P�b%����ËE����   �e���M���e��ËT$�B�J�3��;���H{�]�����������������������������������h(  h��E�P�E�P��$����ËE����   �e���M��me��ËT$�B�J�3��:����z�\�����������������������������������h�   h���E�P�E�P�$����ËE����   �e���M���d��ËT$�B�J�3��4:����{�+\�����������������������������������h�  h���E�P�E�P�$����ËE����   �e���M��d��ËT$�B�J�3���9����}�[����������������������������������̍M��J���T$�B�J�3��9���@}�w[��������������̍������������������M��(���M��w(�������������M��d(��������H ����x����,6����|������   ��|������l����6��Í�T�����5����|������   ��|����������� (��Ë�|������   ��|������������'��Ë�|������   ��|������,����'��Ë�|������   ��|�������'��Í�d����'���M��'��������j����<����N5����|����� �   ��|���ߍ�`����-5��Í�H����!5���T$�B��@���3���7���J�3���7���,w��Y���������������������������������������������������������������������������������������������������������������̋T$�B�J�3��h7���J�3��^7����z�UY������������̋T$�B�J�3��87���L|�/Y����������������������̍M��_���T$�B�J�3�� 7��� ~��X���������������j'h؝�E�P�E�P�� �����j(h؝�E�P�E�P�� �����j)h؝�E�P�E�P�� �����j*h؝�E�P�E�P� �����j+h؝�E�P�E�P� �����j,h؝�E�P�E�P�} �����j-h؝�E�P�E�P�e �����j.h؝��x���P�E�P�J ����ËT$�B��|���3��6���Lt�	X����������������������������������������������������������������̍M�����M�����T$�B�J�3��5��� t�W����������������������̍M����T$�B�J�3��p5����y�gW��������������̍M$�$��������������t��������M��g$���M��_$���M��W$��������*2����$����2��������2���������	2����������1����������1����������1����������1���� �����1���T$�B��t���3��4���J�3��4��� y�V����������������������������������������������������������������̍M��#���T$�B�J�3��@4���J�3��64����v�-V��������������������̍M��E#���T$�B�J�3�� 4���J�3���3���w��U��������������������̍M�����T$�B�J�3���3���}�U��������������̍M��Z���T$�B�J�3��3����|�U��������������̍M��*���T$�B�J�3��`3����|�WU��������������̍M������T$�B�J�3��03����|�'U��������������̍M������M��="���T$�B�J�3���2���J�3���2����x��T����������������������������̍M��z���M���!���T$�B�J�3��2���J�3��2����x�T����������������������������̍M��!���M��{/���T$�B�J�3��X2���J�3��N2���X~�ET����������������������������̍M��U!���M��+/���M��#/���T$�B�J�3�� 2���J�3���1���Xu��S��������������������̍M,��.���M ��.���M�����M�����M�������p����.���M�������|��������d����.���M�����T$�B��l���3��l1����s�cS������������������������������������������̋T$�B�J�3��(1���D��S����������������������̍M��G,���T$�B�J�3���0���`���R��������������̍M��,���T$�B�J�3���0�����R��������������̡��������ËT$�B�J�3��0���P��R������������������������̍M��+���T$�B�J�3��P0������GR��������������̍M��w+���T$�B�J�3�� 0���0��R��������������̍M��G+���T$�B�J�3���/���`���Q�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U����   SVW��@����0   �����������_^[���   ;��8����]���������������������U����   SVW��@����0   ������������_^[���   ;��G8����]���������������������U����   SVW��@����0   ����������L��_^[���   ;���7����]���������������������U����   SVW��@����0   ���������}��_^[���   ;��7����]���������������������U�����L"��]������������������U�����t��]������������������U��������]������������������U�����L��]������������������U�������]������������������U�������]������������������U�����K��]������������������U�칒����]������������������U�친��u���]������������������U�����t��]������������������U��������]������������������U�����K��]������������������U�������]������������������U�������]������������������U�����J��]������������������U�������]������������������U�����"��]������������������U�����MJ��]������������������U�����T��]������������������U��������]������������������U������I��]������������������U��G������]������������������U��D����]������������������U�������]������������������U�����"��]������������������U�����MI��]������������������U�����T��]������������������U��������]������������������U������H��]������������������U��������]������������������U�����b��]������������������U�����H��]������������������U�������]������������������U�������]������������������U�����-H��]��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                            P� ���    ��� ��� � �`�����`�@������� �@����� � ����������0�p�P��0�                                                                                                                                                                                                                                                                                            ������������p�                                                                                                                                                                                                                                                                        `� �    p���0���0��������� ���������    0�p�����    � �    ����    p�`�     ��    0�0���    `�P�    0� �    `�P�    ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �q (T?�D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            c&�$                                                                                                                                                                                                                                                                    ^                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    [ǵZ       s   �
 ��     [ǵZ          �
 �� h74�A�h�06]-9+@<�5        c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ x u t i l i t y                               I T E R A T O R   L I S T   C O R R U P T E D !             �����#�k    bad locale name     p�$�_�_    �@�Ae    c:\program files (x86)\microsoft visual studio 12.0\vc\include\xlocale                  $[j�Ae�&BG*d            c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ x l o c a l e                                 ��.�Ae    �&;�Ae�&7u"0�C3�^.t�Y            H-\�_�_�_�P�&        ��'�k    :    M�k    d1g�F�7�_�P�&        generic     unknown error   ��O�3�n�_�P�&        iostream    iostream stream error        �25O�`rX�P�&        system  ��L�k    d9    ios_base::badbit set        ios_base::failbit set       ios_base::eofbit set            c:\program files (x86)\microsoft visual studio 12.0\vc\include\xiosbase                 ��Q    |�#               $N^-�7] W�A�>k�/g=BeG)[�j�8            Lv6hl�f3Q�>�A�[�!�/g`o�/mX�X�g            �4F        p       ERROR: COULD NOT READ FILE      P�,�)�h�06]-9+@<�5        Load .stl File      STL solid   Ascii stl Files Not Supported!              c:\program files\maxon\cinema 4d r13\plugins\stl_importer\source\stl_importer.cpp                   STL Importer    stl_icon.png        c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ x s t r i n g                                     c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ i s t r e a m                                     c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ v e c t o r                               v e c t o r   s u b s c r i p t   o u t   o f   r a n g e               Standard C++ Libraries Out of Range             " S t a n d a r d   C + +   L i b r a r i e s   O u t   o f   R a n g e "   & &   0                     % s     s t d : : v e c t o r < s t r u c t   t r i a n g l e , c l a s s   s t d : : a l l o c a t o r < s t r u c t   t r i a n g l e >   > : : o p e r a t o r   [ ]                                     " o u t   o f   r a n g e "         ��%�AeD6BG*d�%..mNIJ        i >= 0 && i < count         c:\program files\maxon\cinema 4d r13\resource\_api\ge_dynamicarray.h                %s(%d): %s      string too long     invalid string position         c:\program files (x86)\microsoft visual studio 12.0\vc\include\streambuf                vector<T> too long      s t r i n g   i t e r a t o r   n o t   d e r e f e r e n c a b l e                     s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < c h a r >   >   > : : o p e r a t o r   *                                             i n v a l i d   n u l l   p o i n t e r             bad cast    i n v a l i d   i t e r a t o r   r a n g e             FALSE   c : \ p r o g r a m   f i l e s   ( x 8 6 ) \ m i c r o s o f t   v i s u a l   s t u d i o   1 2 . 0 \ v c \ i n c l u d e \ x m e m o r y                                                           �?        c:\program files\maxon\cinema 4d r13\resource\_api\c4d_resource.cpp                 #   M_EDITOR        c:\program files\maxon\cinema 4d r13\resource\_api\c4d_memory.cpp               c:\program files\maxon\cinema 4d r13\resource\_api\c4d_general.h                   %s  c:\program files\maxon\cinema 4d r13\resource\_api\c4d_string.cpp               no baselist      GB  MB  KB  B        �@    �9i    c:\program files\maxon\cinema 4d r13\resource\_api\c4d_file.cpp             res       �?    ��Mt     �_    x*n        c:\program files\maxon\cinema 4d r13\resource\_api\c4d_baseobject.cpp               nncnt<ncnt      nncnt==ncnt         ����MbP?        c:\program files\maxon\cinema 4d r13\resource\_api\c4d_pmain.cpp                c:\program files\maxon\cinema 4d r13\resource\_api\c4d_basebitmap.cpp               c:\program files\maxon\cinema 4d r13\resource\_api\ge_sort.cpp              c:\program files\maxon\cinema 4d r13\resource\_api\c4d_libs\lib_ngon.cpp                ������        �������    �0m    ,�i    ��U    c:\program files\maxon\cinema 4d r13\resource\_api\c4d_gv\ge_mtools.cpp                 ��i                                                                                                         	           	         	       �d     �d     �d   H   �d       �d      �d      �d     �d      �d   �  e      e   H   e   H   e       e   ��  $e   �                                                           	   alnum   alpha   blank   cntrl   d   digit   graph   lower   print   punct   space  s   upper   w   xdigit  ?          @      @f     Pf     df   H   tf       �f      �f      �f     �f      �f   �  �f      �f   H   �f   H   �f      �f   ��   g   �                                                             	   �   &   ����a l n u m       a l p h a       ����b l a n k       c n t r l       d   d i g i t       g r a p h       l o w e r       p r i n t       p u n c t       s p a c e       s   u p p e r       w   x d i g i t     5            4  �������5            4  �������                   @   �                           0   @   �  �      0                                 @   �                                                        ?                                                                            8�q�k    bad allocation      ��k�k    ��'�k    P�Z�k    �qO�k    �D�k    p�7�c    bad function call       ��s�k        regex_error(error_collate): The expression contained an invalid collating element name.                         regex_error(error_ctype): The expression contained an invalid character class name.                     regex_error(error_escape): The expression contained an invalid escaped character, or a trailing escape.                         regex_error(error_backref): The expression contained an invalid back reference.                 regex_error(error_brack): The expression contained mismatched [ and ].                  regex_error(error_paren): The expression contained mismatched ( and ).                  regex_error(error_brace): The expression contained mismatched { and }.                  regex_error(error_badbrace): The expression contained an invalid range in a { expression }.                     regex_error(error_range): The expression contained an invalid character range, such as [b-a] in most encodings.                         regex_error(error_space): There was insufficient memory to convert the expression into a finite state machine.                          regex_error(error_badrepeat): One of *?+{ was not preceded by a valid regular expression.                       regex_error(error_complexity): The complexity of an attempted match against a regular expression exceeded a pre-set level.                              regex_error(error_stack): There was insufficient memory to determine whether the regular expression could match the specified character sequence.                               regex_error(error_parse)        regex_error(error_syntax)       regex_error     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x s t r i n g                   f:\dd\vctools\crt\crtw32\stdcpp\_tolower.c          f:\dd\vctools\crt\crtw32\stdcpp\locale0.cpp         ,du�Ae    *   C   f:\dd\vctools\crt\crtw32\stdhpp\xutility                      @v�   Xv   hvo   |v�   �v�   �vR   @v�  �v�  �v�  �v   @v7   hvd	  �v�   �v  �vp   �vP   Xv    w'   �v   @v   hv    w   �v{   �v!   <w�   <w�   �v�  @v   Tw   lw   �wn   �va	  �v�  �w   Tw    w   �v�  lw   �v    @v   �w   �v   @v'  �w@'  �wA'  x?'  $x5'  Hx'  pxE'  �xM'  �xF'  �x7'  �x'  �xQ'   y4'  y'  0y&'  @yH'  Ty('  ly8'  �yO'  �yB'  �yD'  �yC'  �yG'  �y:'  �yI'  z6'   z='  0z;'  Lz9'  hzL'  �z3'  �z        f   �zd   �ze   �zq   �z   {!   0{   L{	   \{h   t{    �{j   �{g   �{k   �{l   �{   �wm    |   �v)   �v   $|   Xv   @|&   |v(    wn   T|o   h|*   �|   �|   0y   �v   �|   �v   �|s   �|t   �|u   }v   }w   4}
   H}y   \}'   <wx   h}z   �}{   �}   �v|   �}   �}   hv    w   �}   �}�   ~}   ~~   ,~   Tw�   <~i   �wp   L~   h~�   �~�   �~�   �~   @v�   �~�   �~   �~$      lw"   <   T�   p�   ��   �   �   �w   �r   ��    ��   �                                                                                                                                                                                                                                                                permission denied       file exists     no such device      filename too long       device or resource busy     io error    directory not empty     invalid argument    no space on device      no such file or directory       function not supported      no lock available       not enough memory       resource unavailable try again          cross device link       operation canceled      too many files open     permission_denied       address_in_use      address_not_available       address_family_not_supported        connection_already_in_progress          bad_file_descriptor     connection_aborted      connection_refused      connection_reset    destination_address_required        bad_address     host_unreachable    operation_in_progress       interrupted     invalid_argument    already_connected       too_many_files_open     message_size    filename_too_long       network_down    network_reset   network_unreachable     no_buffer_space     no_protocol_option      not_connected   not_a_socket    operation_not_supported     protocol_not_supported      wrong_protocol_type     timed_out   operation_would_block       address family not supported        address in use      address not available       already connected       argument list too long      argument out of domain      bad address     bad file descriptor     bad message     broken pipe     connection aborted      connection already in progress          connection refused      connection reset    destination address required        executable format error     file too large      host unreachable    identifier removed      illegal byte sequence       inappropriate io control operation          invalid seek    is a directory      message size    network down    network reset   network unreachable     no buffer space     no child process    no link     no message available        no message      no protocol option      no stream resources     no such device or address       no such process     not a directory     not a socket    not a stream    not connected   not supported   operation in progress       operation not permitted     operation not supported     operation would block       owner dead      protocol error      protocol not supported      read only file system       resource deadlock would occur       result out of range     state not recoverable       stream timeout      text file busy      timed out   too many files open in system       too many links      too many symbolic link levels       value too large     wrong protocol type         ��������                    �� e e����������������������                r   a   rb  wb  ab  r+  w+  a+  r+b w+b a+b ��f�f����$�,�4�<�D�P�\�                r   a   r b     w b     a b     r +     w +     a +     r + b       w + b       a + b                
   !   "   2   *            #   3   +                            
   !   "   2   *            #   3   +                   false   true    f:\dd\vctools\crt\crtw32\stdhpp\xlocale         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x l o c a l e                   f:\dd\vctools\crt\crtw32\stdhpp\xlocnum         f:\dd\vctools\crt\crtw32\stdcpp\locale.cpp          �v@�Ae�&�)�(�(�.�.)V)[)�(e.            �n�Ae�C�()�a�a�(�(Ka            Lj�AelO�nskE]{^            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x l o c n u m                   ld  lu  Ld  Lu  %p  0123456789ABCDEFabcdef-+Xx      0123456789-+Ee      eE  pP  .   s t r i n g   s u b s c r i p t   o u t   o f   r a n g e               0123456789ABCDEFabcdef-+XxPp        f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ s t r e a m b u f                       i s t r e a m b u f _ i t e r a t o r   i s   n o t   d e r e f e r e n c a b l e                       i s t r e a m b u f _ i t e r a t o r   i s   n o t   i n c r e m e n t a b l e                         z�����8            _�B        �M�raB3G        f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x u t i l i t y                         :Sun:Sunday:Mon:Monday:Tue:Tuesday:Wed:Wednesday:Thu:Thursday:Fri:Friday:Sat:Saturday                   :Jan:January:Feb:February:Mar:March:Apr:April:May:May:Jun:June:Jul:July:Aug:August:Sep:September:Oct:October:Nov:November:Dec:December                                  : S u n : S u n d a y : M o n : M o n d a y : T u e : T u e s d a y : W e d : W e d n e s d a y : T h u : T h u r s d a y : F r i : F r i d a y : S a t : S a t u r d a y                                       : J a n : J a n u a r y : F e b : F e b r u a r y : M a r : M a r c h : A p r : A p r i l : M a y : M a y : J u n : J u n e : J u l : J u l y : A u g : A u g u s t : S e p : S e p t e m b e r : O c t : O c t o b e r : N o v : N o v e m b e r : D e c : D e c e m b e r                                                         �pZ�Ae�(!6,+�]�H�6|N        �!�AeS�Q�(�l�]M(#C        ti%�AeXY0,3�u�L4Z�^pd5r�.�a�Q            �|]�Aeud�$R_^:�joL�%'�$�a(1D            ����\�H�Ae    ��+�Ae     �i�Ae    �#�=�Ae�Y    f:\dd\vctools\crt\crtw32\stdcpp\wlocale.cpp         <7>�Ae�g)j�i�i�%8$-kej2k~j&            | 8�Ae�+\ \�4�4�Y*Z�4            ��>�Ae4<�i d�E�T        � �+�Aes�n
f        <!(k�Aenf@�         �!�R�Ae�5�X     "�Q�Ae�a�]    H$�E�Ae?J�<;q�27%�0 MsH�;            `"Hs�Ae?J�<;q�27%�0 MsH�;            #A9�Ae?J�<;q�27%�0 MsH�;            �#fn�Ae�Ex96ObB�]+6        �3L�Ae�%!'&'�&[[[#%(%%Z%V[            `$6q�Ae'u2�2NrDr�2�2�q            �$56�Ae�'�>�[;+�*         %�k�Ae�:�A�s        �%.=�Ae�8mDR-        �%\-�Aec5�;    ����D&%2�AeSEc0    �(k#�AeVtdH@g�5�d�406�(�"            �&SY�AeVtdH@g�5�d�406�(�"            \'yG�AeVtdH@g�5�d�406�(�"            �'K�Ae,�_o�5P4FC�>        ,(�;�AexR    f:\dd\vctools\crt\crtw32\stdhpp\xloctime            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x l o c t i m e                     ! % x       f:\dd\vctools\crt\crtw32\stdhpp\locale          f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ l o c a l e                     f:\dd\vctools\crt\crtw32\stdhpp\xlocmes         f:\dd\vctools\crt\crtw32\stdhpp\xlocmon         %.0Lf   0123456789-     %b %d %H : %M : %S %Y       %m / %d / %y        :AM:am:PM:pm    %I : %M : %S %p     %H : %M     %H : %M : S     %d / %m / %y    0123456789-     0123456789ABCDEFabcdef-+Xx      0123456789-+Ee          f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d h p p \ x l o c m o n                   0123456789-     0123456789ABCDEFabcdef-+Xx      0123456789-+Ee      0123456789-     0123456789ABCDEFabcdef-+XxPp        $+xv    : A M : a m : P M : p m         0123456789ABCDEFabcdef-+XxPp            s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < w c h a r _ t >   >   > : : o p e r a t o r   *                                               s t r i n g   i t e r a t o r   n o t   i n c r e m e n t a b l e                       s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < w c h a r _ t >   >   > : : o p e r a t o r   + +                                             s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < u n s i g n e d   s h o r t >   >   > : : o p e r a t o r   *                                                 s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < u n s i g n e d   s h o r t >   >   > : : o p e r a t o r   + +                                                   -   +v$x+v$xv$+xv+$xv$+x+$vx+$vx$v+x+$vx$+vx+v $+v $v $+v +$v $++$ v+$ v$ v++$ v$+ v+xv$+ v$v$ +v+ $v$ ++x$v+ $v$v ++ $v$ +v                                s t r i n g   i t e r a t o r   +   o f f s e t   o u t   o f   r a n g e                       s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < w c h a r _ t >   >   > : : o p e r a t o r   + =                                             s t r i n g   i t e r a t o r s   i n c o m p a t i b l e               Standard C++ Libraries Invalid Argument         " S t a n d a r d   C + +   L i b r a r i e s   I n v a l i d   A r g u m e n t "   & &   0                     s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < w c h a r _ t >   >   > : : _ C o m p a t                                             " i n v a l i d   a r g u m e n t "             s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < u n s i g n e d   s h o r t >   >   > : : o p e r a t o r   + =                                               s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < u n s i g n e d   s h o r t >   >   > : : _ C o m p a t                                               -   �(�M�Ae%�r�i        f:\dd\vctools\crt\crtw32\stdcpp\xlocale.cpp         )pP�Ae�O|bPC        h),D�Ae�n�H    �)�A�Ae�@}%    ,_C�AeW�n�S�P�f�d>�5�N            (*{c�AeW�n�S�P�f�d>�5�N            �*�F�AeW�n�S�P�f�d>�5�N            L+J:�Aeje�$Vov,	IZ/P         �+;5�Ae.)    0123456789-     !%x     0123456789-         s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < c h a r >   >   > : : o p e r a t o r   + +                                           s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < c h a r >   >   > : : o p e r a t o r   + =                                           s t d : : _ S t r i n g _ c o n s t _ i t e r a t o r < c l a s s   s t d : : _ S t r i n g _ v a l < s t r u c t   s t d : : _ S i m p l e _ t y p e s < c h a r >   >   > : : _ C o m p a t                                                 �M(knN          �A            e��A    0123456789abcdefghijklmnopqrstuvwxyz      !

					               0123456789abcdefghijklmnopqrstuvwxyz      A)!                   p l o c - > _ M b c u r m a x   = =   1   | |   p l o c - > _ M b c u r m a x   = =   2                         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d c p p \ x m b t o w c . c                   f:\dd\vctools\crt\crtw32\stdcpp\xwcsxfrm.c          0123456789abcdefABCDEF   	

            �?  �? @F   �  �� ��= �9 �3       A      �?              �              �           ����?   ���9>   033�<              $@           ����?   ���9>   033�<           ?  � ������?�                      ?  � ������?�                         f:\dd\vctools\crt\crtw32\misc\onexit.c          ����    d s t   ! =   N U L L       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ m e m c p y _ s . c                     m e m c p y _ s         s r c   ! =   N U L L       s i z e I n B y t e s   > =   c o u n t             (,A/�k    Unknown exception       @,�,�k    �,H�k    �,�p�k    ( s t r e a m   ! =   N U L L )         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f c l o s e . c                   f c l o s e     ( s t r   ! =   N U L L )           _ f c l o s e _ n o l o c k         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f g e t c . c                     f g e t c       (   ( _ S t r e a m - > _ f l a g   &   _ I O S T R G )   | |   (   f n   =   _ f i l e n o ( _ S t r e a m ) ,   (   ( _ t e x t m o d e _ s a f e ( f n )   = =   _ _ I O I N F O _ T M _ A N S I )   & &   ! _ t m _ u n i c o d e _ s a f e ( f n ) ) ) )                                                       g e t c     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f g e t p o s . c                     f g e t p o s       ( p o s   ! =   N U L L )               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f p u t c . c                     f p u t c       p u t c         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f s e t p o s . c                     f s e t p o s       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f s e e k i 6 4 . c                   _ f s e e k i 6 4           ( ( w h e n c e   = =   S E E K _ S E T )   | |   ( w h e n c e   = =   S E E K _ C U R )   | |   ( w h e n c e   = =   S E E K _ E N D ) )                                 s t r   ! =   N U L L       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f w r i t e . c                   f w r i t e     _ f w r i t e _ n o l o c k         ( b u f f e r   ! =   N U L L )         n u m   < =   ( S I Z E _ M A X   /   s i z e )             ( " I n c o n s i s t e n t   S t r e a m   C o u n t .   F l u s h   b e t w e e n   c o n s e c u t i v e   r e a d   a n d   w r i t e " ,   s t r e a m - > _ c n t   > =   0 )                                             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ s e t v b u f . c                     s e t v b u f       ( t y p e   = =   _ I O N B F )   | |   ( t y p e   = =   _ I O F B F )   | |   ( t y p e   = =   _ I O L B F )                         ( ( 2   < =   s i z e )   & &   ( s i z e   < =   I N T _ M A X ) )                 f:\dd\vctools\crt\crtw32\stdio\setvbuf.c            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ u n g e t c . c                   u n g e t c     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ u n g e t c _ n o l o c k . i n l                     _ u n g e t c _ n o l o c k         f:\dd\vctools\crt\crtw32\stdio\_file.c          0�D�T�    W a r n i n g       E r r o r       A s s e r t i o n   F a i l e d         . . .       m o d e   = =   _ C R T _ R P T H O O K _ I N S T A L L   | |   m o d e   = =   _ C R T _ R P T H O O K _ R E M O V E                           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ d b g r p t . c                     _ C r t S e t R e p o r t H o o k W 2           p f n N e w H o o k   ! =   N U L L             ( " T h e   h o o k   f u n c t i o n   i s   n o t   i n   t h e   l i s t ! " , 0 )                       f:\dd\vctools\crt\crtw32\misc\dbgrpt.c          _ _ c r t M e s s a g e W i n d o w W               w c s c p y _ s ( s z E x e N a m e ,   2 6 0 ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                       < p r o g r a m   n a m e   u n k n o w n >                 m e m c p y _ s ( s z S h o r t P r o g N a m e ,   s i z e o f ( T C H A R )   *   ( 2 6 0   -   ( s z S h o r t P r o g N a m e   -   s z E x e N a m e ) ) ,   d o t d o t d o t ,   s i z e o f ( T C H A R )   *   3 )                                                     
 
 F o r   i n f o r m a t i o n   o n   h o w   y o u r   p r o g r a m   c a n   c a u s e   a n   a s s e r t i o n 
 f a i l u r e ,   s e e   t h e   V i s u a l   C + +   d o c u m e n t a t i o n   o n   a s s e r t s .                                                 E x p r e s s i o n :           
 
     
 L i n e :         
 F i l e :         
 M o d u l e :             D e b u g   % s ! 
 
 P r o g r a m :   % s % s % s % s % s % s % s % s % s % s % s % s 
 
 ( P r e s s   R e t r y   t o   d e b u g   t h e   a p p l i c a t i o n ) 
                                       ( * _ e r r n o ( ) )           w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r                     M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y                 p�x�������    Free    Normal  CRT Ignore  Client  _ C r t C h e c k M e m o r y ( )           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ d b g h e a p . c                   Client hook allocation failure at file %hs line %d.
            Client hook allocation failure.
        Invalid allocation size: %Iu bytes.
        Error: memory allocation: bad memory block type.
           Client hook re-allocation failure at file %hs line %d.
             Client hook re-allocation failure.
         Invalid allocation size: %Iu bytes.

Memory allocated at %hs(%d).
              Error: memory allocation: bad memory block type.

Memory allocated at %hs(%d).
                 The Block at 0x%p was allocated by aligned routines, use _aligned_realloc()                     _ C r t I s V a l i d H e a p P o i n t e r ( p U s e r D a t a )                       p O l d B l o c k - > n L i n e   = =   I G N O R E _ L I N E   & &   p O l d B l o c k - > l R e q u e s t   = =   I G N O R E _ R E Q                                 Error: possible heap corruption at or near 0x%p                 f R e a l l o c   | |   ( ! f R e a l l o c   & &   p N e w B l o c k   = =   p O l d B l o c k )                       _ p L a s t B l o c k   = =   p O l d B l o c k             _ p F i r s t B l o c k   = =   p O l d B l o c k               p U s e r D a t a   ! =   N U L L           _ e x p a n d _ d b g           The Block at 0x%p was allocated by aligned routines, use _aligned_free()                Client hook free failure.
      _ B L O C K _ T Y P E _ I S _ V A L I D ( p H e a d - > n B l o c k U s e )                     HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.

Memory allocated at %hs(%d).
                                         HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.
                               HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.

Memory allocated at %hs(%d).
                                     HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.
                           p H e a d - > n L i n e   = =   I G N O R E _ L I N E   & &   p H e a d - > l R e q u e s t   = =   I G N O R E _ R E Q                             p H e a d - > n B l o c k U s e   = =   n B l o c k U s e               _ p L a s t B l o c k   = =   p H e a d             _ p F i r s t B l o c k   = =   p H e a d           _ m s i z e _ d b g         _heapchk fails with _HEAPBADBEGIN.
         _heapchk fails with _HEAPBADNODE.
          _heapchk fails with _HEAPBADEND.
       _heapchk fails with _HEAPBADPTR.
       _heapchk fails with unknown return value!
          DAMAGED     HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.

Memory allocated at %hs(%d).
                                 HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.
                               %hs located at 0x%p is %Iu bytes long.

Memory allocated at %hs(%d).
               %hs located at 0x%p is %Iu bytes long.
             ( f N e w B i t s = = _ C R T D B G _ R E P O R T _ F L A G )   | |   ( ( f N e w B i t s   &   0 x 0 f f f f   &   ~ ( _ C R T D B G _ A L L O C _ M E M _ D F   |   _ C R T D B G _ D E L A Y _ F R E E _ M E M _ D F   |   _ C R T D B G _ C H E C K _ A L W A Y S _ D F   |   _ C R T D B G _ C H E C K _ C R T _ D F   |   _ C R T D B G _ L E A K _ C H E C K _ D F )   )   = =   0 )                                                                                 _ C r t S e t D b g F l a g         p f n   ! =   N U L L       _ C r t D o F o r A l l C l i e n t O b j e c t s               s t a t e   ! =   N U L L           _ C r t M e m C h e c k p o i n t           Bad memory block found at 0x%p.

Memory allocated at %hs(%d).
              Bad memory block found at 0x%p.
        _ C r t M e m D i f f e r e n c e           o l d S t a t e   ! =   N U L L         n e w S t a t e   ! =   N U L L         %.2X    _ p r i n t M e m B l o c k D a t a              Data: <%s> %s
     Dumping objects ->
     #File Error#(%d) :      %hs(%d) :       {%ld}   client block at 0x%p, subtype %x, %Iu bytes long.
              normal block at 0x%p, %Iu bytes long.
          crt block at 0x%p, subtype %x, %Iu bytes long.
             Object dump complete.
      Detected memory leaks!
     _ C r t M e m D u m p S t a t i s t i c s           %Id bytes in %Id %hs Blocks.
       Largest number used: %Id bytes.
        Total allocations: %Id bytes.
          I S _ 2 _ P O W _ N ( a l i g n )           _ a l i g n e d _ o f f s e t _ m a l l o c _ d b g             o f f s e t   = =   0   | |   o f f s e t   <   s i z e                 The block at 0x%p was not allocated by _aligned routines, use realloc()                 Damage before 0x%p which was allocated by aligned routine
              _ a l i g n e d _ o f f s e t _ r e a l l o c _ d b g                   The block at 0x%p was not allocated by _aligned routines, use free()                m e m b l o c k   ! =   N U L L         _ a l i g n e d _ m s i z e _ d b g             csm�               �                X- R    �S    f:\dd\vctools\crt\crtw32\startup\dllcrt0.c                            �A������               �             ��      �C      �C   ����G   ���8      `E           � 3  ?     �  ?                          f:\dd\vctools\crt\crtw32\startup\mlock.c            ;�-1X�k    bad exception                                                                                                                                                                                                                                                                                         ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               ( ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                                                            �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ w c s d u p . c                     _ w c s d u p _ d b g       w c s c p y _ s ( m e m o r y ,   s i z e ,   s t r i n g )                 f:\dd\vctools\crt\crtw32\misc\initctyp.c            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ i n i t c t y p . c                     p l o c i - > c t y p e 1 _ r e f c o u n t   >   0                 ( " C o r r u p t e d   p o i n t e r   p a s s e d   t o   _ f r e e a " ,   0 )                       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ m a l l o c . h                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ s e t l o c a l . c                     s e t l o c a l e           m b s t o w c s _ s ( & s i z e ,   ( ( v o i d   * ) 0 ) ,   0 ,   _ l o c a l e ,   2 1 4 7 4 8 3 6 4 7 )                         f:\dd\vctools\crt\crtw32\misc\setlocal.c            m b s t o w c s _ s ( ( ( v o i d   * ) 0 ) ,   i n w l o c a l e ,   s i z e ,   _ l o c a l e ,   ( ( s i z e _ t ) - 1 ) )                                   _ w c s t o m b s _ s _ l ( & s i z e ,   ( ( v o i d   * ) 0 ) ,   0 ,   o u t w l o c a l e ,   0 ,   & l o c a l e )                                 _ w c s t o m b s _ s _ l ( ( ( v o i d   * ) 0 ) ,   o u t l o c a l e ,   s i z e ,   o u t w l o c a l e ,   ( ( s i z e _ t ) - 1 ) ,   & l o c a l e )                                     ( ( p t l o c i - > l c _ c a t e g o r y [ _ c a t e g o r y ] . l o c a l e   ! =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ _ c a t e g o r y ] . r e f c o u n t   ! =   N U L L ) )   | |   ( ( p t l o c i - > l c _ c a t e g o r y [ _ c a t e g o r y ] . l o c a l e   = =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ _ c a t e g o r y ] . r e f c o u n t   = =   N U L L ) )                                                                                         ( f i l e   ! =   N U L L )             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f o p e n . c                     _ f s o p e n       ( m o d e   ! =   N U L L )         ( * m o d e   ! =   _ T ( ' \ 0 ' ) )           ( p f i l e   ! =   N U L L )           f o p e n _ s           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f s e e k . c                     f s e e k       _ w f s o p e n         _ w f o p e n _ s       k e r n e l 3 2 . d l l         FlsAlloc    FlsFree     FlsGetValue     FlsSetValue     InitializeCriticalSectionEx         CreateEventExW      CreateSemaphoreExW      SetThreadStackGuarantee     CreateThreadpoolTimer       SetThreadpoolTimer      WaitForThreadpoolTimerCallbacks         CloseThreadpoolTimer        CreateThreadpoolWait        SetThreadpoolWait       CloseThreadpoolWait     FlushProcessWriteBuffers        FreeLibraryWhenCallbackReturns          GetCurrentProcessorNumber       GetLogicalProcessorInformation          CreateSymbolicLinkW     SetDefaultDllDirectories        EnumSystemLocalesEx     CompareStringEx     GetDateFormatEx     GetLocaleInfoEx     GetTimeFormatEx     GetUserDefaultLocaleName        IsValidLocaleName       LCMapStringEx   GetCurrentPackageId     GetTickCount64      GetFileInformationByHandleExW       SetFileInformationByHandleW         ( f o r m a t   ! =   N U L L )             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ s p r i n t f . c                     s p r i n t f       ( s t r i n g   ! =   N U L L )         p V a l u e   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ d o s \ d o s m a p . c                   _ g e t _ e r r n o         _ g e t _ d o s e r r n o           f:\dd\vctools\crt\crtw32\time\strftime.c            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ t i m e \ s t r f t i m e . c                     _ G e t d a y s _ l         s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > w d a y _ a b b r [ n ] )                             s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > w d a y [ n ] )                       _ G e t m o n t h s _ l         s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > m o n t h _ a b b r [ n ] )                           s t r c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > m o n t h [ n ] )                     (   s t r i n g   ! =   N U L L   )             _ S t r f t i m e _ l       (   m a x s i z e   ! =   0   )         (   f o r m a t   ! =   N U L L   )             (   t i m e p t r   ! =   N U L L   )           f:\dd\vctools\crt\crtw32\time\wcsftime.c            f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ t i m e \ w c s f t i m e . c                     _ W _ G e t d a y s _ l             w c s c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > _ W _ w d a y _ a b b r [ n ] )                               w c s c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > _ W _ w d a y [ n ] )                         _ W _ G e t m o n t h s _ l             w c s c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > _ W _ m o n t h _ a b b r [ n ] )                             w c s c p y _ s ( s ,   ( l e n   +   1 )   -   ( s   -   p ) ,   p t - > _ W _ m o n t h [ n ] )                       _ W _ G e t t n a m e s _ l             s t r c p y _ s ( d e s t - > w d a y _ a b b r [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > w d a y _ a b b r [ i d x ] )                                       s t r c p y _ s ( d e s t - > w d a y [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > w d a y [ i d x ] )                                   s t r c p y _ s ( d e s t - > m o n t h _ a b b r [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > m o n t h _ a b b r [ i d x ] )                                           s t r c p y _ s ( d e s t - > m o n t h [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > m o n t h [ i d x ] )                                       s t r c p y _ s ( d e s t - > a m p m [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > a m p m [ i d x ] )                                   s t r c p y _ s ( d e s t - > w w _ s d a t e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > w w _ s d a t e f m t )                                           s t r c p y _ s ( d e s t - > w w _ l d a t e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > w w _ l d a t e f m t )                                           s t r c p y _ s ( d e s t - > w w _ t i m e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( c h a r ) ,   s r c - > w w _ t i m e f m t )                                       w c s c p y _ s ( d e s t - > _ W _ w d a y _ a b b r [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w d a y _ a b b r [ i d x ] )                                             w c s c p y _ s ( d e s t - > _ W _ w d a y [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w d a y [ i d x ] )                                         w c s c p y _ s ( d e s t - > _ W _ m o n t h _ a b b r [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ m o n t h _ a b b r [ i d x ] )                                                 w c s c p y _ s ( d e s t - > _ W _ m o n t h [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ m o n t h [ i d x ] )                                             w c s c p y _ s ( d e s t - > _ W _ a m p m [ i d x ] ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ a m p m [ i d x ] )                                         w c s c p y _ s ( d e s t - > _ W _ w w _ s d a t e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w w _ s d a t e f m t )                                         w c s c p y _ s ( d e s t - > _ W _ w w _ l d a t e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w w _ l d a t e f m t )                                         w c s c p y _ s ( d e s t - > _ W _ w w _ t i m e f m t ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w w _ t i m e f m t )                                             w c s c p y _ s ( d e s t - > _ W _ w w _ l o c a l e _ n a m e ,   ( t o t a l _ b y t e s   -   b y t e s )   /   s i z e o f ( w c h a r _ t ) ,   s r c - > _ W _ w w _ l o c a l e _ n a m e )                                             _ W c s f t i m e _ l       t i m e p t r   ! =   N U L L           F A L S E           (   (   t i m e p t r - > t m _ w d a y   > = 0   )   & &   (   t i m e p t r - > t m _ w d a y   < =   6   )   )                           _ W _ e x p a n d t i m e           (   (   t i m e p t r - > t m _ m o n   > = 0   )   & &   (   t i m e p t r - > t m _ m o n   < =   1 1   )   )                         (   (   t i m e p t r - > t m _ m d a y   > = 1   )   & &   (   t i m e p t r - > t m _ m d a y   < =   3 1   )   )                             (   (   t i m e p t r - > t m _ h o u r   > = 0   )   & &   (   t i m e p t r - > t m _ h o u r   < =   2 3   )   )                             (   (   t i m e p t r - > t m _ y d a y   > = 0   )   & &   (   t i m e p t r - > t m _ y d a y   < =   3 6 5   )   )                           (   (   t i m e p t r - > t m _ m i n   > = 0   )   & &   (   t i m e p t r - > t m _ m i n   < =   5 9   )   )                         (   (   t i m e p t r - > t m _ s e c   > = 0   )   & &   (   t i m e p t r - > t m _ s e c   < =   5 9   )   )                         (   t i m e p t r - > t m _ y e a r   > = 0   )                 (   t i m e p t r - > t m _ y e a r   > =   - 1 9 0 0   )   & &   (   t i m e p t r - > t m _ y e a r   < =   8 0 9 9   )                               _ m b s t o w c s _ s _ l ( & w n u m ,   * s t r i n g ,   * l e f t ,   ( _ _ t z n a m e ( ) ) [ ( ( t i m e p t r - > t m _ i s d s t ) ? 1 : 0 ) ] ,   ( ( s i z e _ t ) - 1 ) ,   p l o c i n f o )                                               (   " I n v a l i d   f o r m a t   d i r e c t i v e "   ,   0   )                 a m / p m       a / p       c c h C o u n t 1 = = 0   & &   c c h C o u n t 2 = = 1   | |   c c h C o u n t 1 = = 1   & &   c c h C o u n t 2 = = 0                                 f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ a _ c m p . c                   c a     z h - C H S     c s     d a     d e     e l     e n     e s     f i     f r     h e     h u     i s     i t     j a     k o     n l     n o     p l     p t     r o     r u     h r     s k     s q     s v     t h     t r     u r     i d     u k     b e     s l     e t     l v     l t     f a     v i     h y     a z     e u     m k     a f     k a     f o     h i     m s     k k     k y     s w     u z     t t     p a     g u     t a     t e     k n     m r     s a     m n     g l     k o k       s y r       d i v       a r - S A       b g - B G       c a - E S       z h - T W       c s - C Z       d a - D K       d e - D E       e l - G R       e n - U S       f i - F I       f r - F R       h e - I L       h u - H U       i s - I S       i t - I T       j a - J P       k o - K R       n l - N L       n b - N O       p l - P L       p t - B R       r o - R O       r u - R U       h r - H R       s k - S K       s q - A L       s v - S E       t h - T H       t r - T R       u r - P K       i d - I D       u k - U A       b e - B Y       s l - S I       e t - E E       l v - L V       l t - L T       f a - I R       v i - V N       h y - A M       a z - A Z - L a t n         e u - E S       m k - M K       t n - Z A       x h - Z A       z u - Z A       a f - Z A       k a - G E       f o - F O       h i - I N       m t - M T       s e - N O       m s - M Y       k k - K Z       k y - K G       s w - K E       u z - U Z - L a t n         t t - R U       b n - I N       p a - I N       g u - I N       t a - I N       t e - I N       k n - I N       m l - I N       m r - I N       s a - I N       m n - M N       c y - G B       g l - E S       k o k - I N     s y r - S Y     d i v - M V     q u z - B O     n s - Z A       m i - N Z       a r - I Q       z h - C N       d e - C H       e n - G B       e s - M X       f r - B E       i t - C H       n l - B E       n n - N O       p t - P T       s r - S P - L a t n         s v - F I       a z - A Z - C y r l         s e - S E       m s - B N       u z - U Z - C y r l         q u z - E C     a r - E G       z h - H K       d e - A T       e n - A U       e s - E S       f r - C A       s r - S P - C y r l         s e - F I       q u z - P E     a r - L Y       z h - S G       d e - L U       e n - C A       e s - G T       f r - C H       h r - B A       s m j - N O     a r - D Z       z h - M O       d e - L I       e n - N Z       e s - C R       f r - L U       b s - B A - L a t n         s m j - S E     a r - M A       e n - I E       e s - P A       f r - M C       s r - B A - L a t n         s m a - N O     a r - T N       e n - Z A       e s - D O       s r - B A - C y r l         s m a - S E     a r - O M       e n - J M       e s - V E       s m s - F I     a r - Y E       e n - C B       e s - C O       s m n - F I     a r - S Y       e n - B Z       e s - P E       a r - J O       e n - T T       e s - A R       a r - L B       e n - Z W       e s - E C       a r - K W       e n - P H       e s - C L       a r - A E       e s - U Y       a r - B H       e s - P Y       a r - Q A       e s - B O       e s - S V       e s - H N       e s - N I       e s - P R       z h - C H T     s r         ��B   $,   t"q   �,    �"�   �"�   �"�   �"�   �"�   �"�   �"�   �"�   #�   #�   $#�   4#�   D#C   T#�   d#�   t#�   )   �#�   �#k   �!   �#c   �,   �#D   �#}   �#�   �   $E   �   $G   ($�   �   8$H   �   H$�   X$�   h$I   x$�   �$�   �A   �$�   �   �$J      �$�   �$�   �$�   �$�   �$�   %�   %�   (%�   8%�   H%�   X%K   h%�   x%�   	   �%�   �%�   �%�   �%�   �%�   �%�   �%�   �%�   &�   &�   (&�   8&�   H&�   X&�   h&�   x&�   �&�   �&�   �&�   �#   �&e   *   �&l   �&   �&h   
   �&L   4.   �&s      '�   '�   ('�   8'M   H'�   X'�   �>   h'�   |7   x'   $   �'N   </   �'t   �   �'�   �'Z   ,   �'O   (   �'j   �   �'a   4   �'P   <   (�   (Q   D   ((R   ,-   8(r   L1   H(x   �:   X(�   L   �?   h(�   x(S   T2   �(y   �%   �(g   �$   �(f   �(�   +   �(m   �(�   �=   �(�   �;   �(�   D0   )�   )w   ()u   8)U   T   H)�   X)T   h)�   \   x)�   t6   �)~   d   �)V   l   �)W   �)�   �)�   �)�   �)�   t   �)X   |   *Y   �<   *�   (*�   8*v   H*�   �   X*[   �"   h*d   x*�   �*�   �*�   �*�   �*�   �*�   �   �*\   L�   �*�   +�    +�   <+�   �   X+�   h+]   \3   x+z   �@   �+�   �8   �+�   �9   �+�   �   �+^   �+n   �   �+_   l5   �+|   �    �+b   �   ,`   d4   ,�   4,{   �'   P,i   `,o   p,   �,�   �,�   �,�   �,�   �,�   �,F   �,p      �,   �,   �   �   �   �   �   �	   
            $   ,   4   <   D   L   T   \   d   l   t   |   �   �   �   �   �   �    �!   �"   �#   �$   �%   �&   �'   �)   �*   �+   ,   -   /   6   $7   ,8   49   <>   D?   L@   TA   \C   dD   lF   tG   |I   �J   �K   �N   �O   �P   �V   �W   �Z   �e   �   ��  �  �          0  @  P	  `  p  �  �  �  �  �  �  �  �          0  @  P  `  p  �  �  �   �!  �"  �#  �$  �%   	&  	'   	)  0	*  @	+  P	,  `	-  |	/  �	2  �	4  �	5  �	6  �	7  �	8  �	9  �	:  
;  
>  ,
?  <
@  L
A  \
C  l
D  �
E  �
F  �
G  �
I  �
J  �
K  �
L  �
N  O  P  (R  8V  HW  XZ  he  xk  �l  ��  �  �  �  �	  �
  �      (  8  H  X  t,  �;  �>  �C  �k  �  �  �  	  
  ,  <  L;  hk  x  �  �  �	  �
  �  �  �;  �      (	  8
  H  X  h;  �  �	  �
  �  �  �;  �   	  
     0;  L   \	   l
   |;   �$  �	$  �
$  �;$  �(  �	(  �
(  �,  	,  
,  ,0  <	0  L
0  \4  l	4  |
4  �8  �
8  �<  �
<  �@  �
@  �
D  �
H  
L  
P  ,|  <|  L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            a f - z a       a r - a e       a r - b h       a r - d z       a r - e g       a r - i q       a r - j o       a r - k w       a r - l b       a r - l y       a r - m a       a r - o m       a r - q a       a r - s a       a r - s y       a r - t n       a r - y e       a z - a z - c y r l         a z - a z - l a t n         b e - b y       b g - b g       b n - i n       b s - b a - l a t n         c a - e s       c s - c z       c y - g b       d a - d k       d e - a t       d e - c h       d e - d e       d e - l i       d e - l u       d i v - m v     e l - g r       e n - a u       e n - b z       e n - c a       e n - c b       e n - g b       e n - i e       e n - j m       e n - n z       e n - p h       e n - t t       e n - u s       e n - z a       e n - z w       e s - a r       e s - b o       e s - c l       e s - c o       e s - c r       e s - d o       e s - e c       e s - e s       e s - g t       e s - h n       e s - m x       e s - n i       e s - p a       e s - p e       e s - p r       e s - p y       e s - s v       e s - u y       e s - v e       e t - e e       e u - e s       f a - i r       f i - f i       f o - f o       f r - b e       f r - c a       f r - c h       f r - f r       f r - l u       f r - m c       g l - e s       g u - i n       h e - i l       h i - i n       h r - b a       h r - h r       h u - h u       h y - a m       i d - i d       i s - i s       i t - c h       i t - i t       j a - j p       k a - g e       k k - k z       k n - i n       k o k - i n     k o - k r       k y - k g       l t - l t       l v - l v       m i - n z       m k - m k       m l - i n       m n - m n       m r - i n       m s - b n       m s - m y       m t - m t       n b - n o       n l - b e       n l - n l       n n - n o       n s - z a       p a - i n       p l - p l       p t - b r       p t - p t       q u z - b o     q u z - e c     q u z - p e     r o - r o       r u - r u       s a - i n       s e - f i       s e - n o       s e - s e       s k - s k       s l - s i       s m a - n o     s m a - s e     s m j - n o     s m j - s e     s m n - f i     s m s - f i     s q - a l       s r - b a - c y r l         s r - b a - l a t n         s r - s p - c y r l         s r - s p - l a t n         s v - f i       s v - s e       s w - k e       s y r - s y     t a - i n       t e - i n       t h - t h       t n - z a       t r - t r       t t - r u       u k - u a       u r - p k       u z - u z - c y r l         u z - u z - l a t n         v i - v n       x h - z a       z h - c h s     z h - c h t     z h - c n       z h - h k       z h - m o       z h - s g       z h - t w       z u - z a       a r     b g     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ w i n a p i n l s . c                   _ _ c r t D o w n l e v e l L C I D T o L o c a l e N a m e                 w c s c p y _ s ( o u t L o c a l e N a m e ,   c c h L o c a l e N a m e ,   b u f f e r )                     �.�/H1l1�1�1                   Stack around the variable ' ' was corrupted.    The variable '  ' is being used without being initialized.                                      The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.
                                                    A cast to a smaller data type has caused a loss of data.  If this was intentional, you should mask the source of the cast with the appropriate bitmask.  For example:  
	char c = (i & 0xFF);
Changing the code in this way will not affect the quality of the resulting optimized code.
                                                            Stack memory was corrupted
        A local variable was used before it was initialized
           Stack memory around _alloca was corrupted
         Unknown Runtime Check Error
           R u n t i m e   C h e c k   E r r o r . 
    U n a b l e   t o   d i s p l a y   R T C   M e s s a g e .                               R u n - T i m e   C h e c k   F a i l u r e   # % d   -   % s               Unknown Filename    Unknown Module Name     Run-Time Check Failure #%d - %s         Stack corrupted near unknown variable           u s e r 3 2 . d l l         wsprintfA   Stack area around _alloca memory reserved by this function is corrupted
                
Data: <    
Allocation number within this function:            
Size:      
Address: 0x        Stack area around _alloca memory reserved by this function is corrupted                 %s%s%p%s%ld%s%d%s       
   >   %s%s%s%s    A variable is being used without being initialized.             5<5p5�5�5    Stack pointer corruption        Cast to smaller type causing loss of data           Stack memory corruption     Local variable used before initialization           Stack around _alloca corrupted          The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.                                              f:\dd\vctools\crt\crtw32\misc\i386\chkesp.c                8   x8	   �8
   P9   �9   :   �:   �:   @;   �;    <   �<    =   x=   �=    �>!   8?"   �Ax   By   (Bz   HB�   lB�   tB                                        R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
                         R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
                       R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
                           R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
                     R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
                           R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
                         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
                 R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
                         R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
                         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
                       R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
                         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
                         R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
                 R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
                     R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
                                             R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
                             R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
                                                                                                     R 6 0 3 4  
 -   i n c o n s i s t e n t   o n e x i t   b e g i n - e n d   v a r i a b l e s  
                         D O M A I N   e r r o r  
         S I N G   e r r o r  
         T L O S S   e r r o r  
            
     r u n t i m e   e r r o r           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t a r t u p \ c r t 0 m s g . c                     _ N M S G _ W R I T E           w c s c p y _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " R u n t i m e   E r r o r ! \ n \ n P r o g r a m :   " )                                     R u n t i m e   E r r o r ! 
 
 P r o g r a m :                 w c s c p y _ s ( p r o g n a m e ,   p r o g n a m e _ s i z e ,   L " < p r o g r a m   n a m e   u n k n o w n > " )                                 w c s n c p y _ s ( p c h ,   p r o g n a m e _ s i z e   -   ( p c h   -   p r o g n a m e ) ,   L " . . . " ,   3 )                           w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " \ n \ n " )                                   w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   e r r o r _ t e x t )                             f:\dd\vctools\crt\crtw32\misc\inithelp.c                f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ i n i t h e l p . c                     _ _ g e t l o c a l e i n f o               s t r n c p y _ s ( * s t r a d d r e s s ,   o u t s i z e ,   p c b u f f e r ,   o u t s i z e   -   1 )                         m s c o r e e . d l l       CorExitProcess          f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t a r t u p \ c r t 0 d a t . c                     _ g e t _ w p g m p t r         _ w p g m p t r   ! =   N U L L         _ g e t _ p g m p t r       _ p g m p t r   ! =   N U L L           p a t h   ! =   N U L L         _ _ c o p y _ p a t h _ t o _ w i d e _ s t r i n g             o u t P a t h   ! =   N U L L           f:\dd\vctools\crt\crtw32\startup\crt0dat.c          i n S t r i n g   ! =   N U L L         _ _ c o p y _ t o _ c h a r         o u t S t r i n g   ! =   N U L L           exp pow log log10   sinh    cosh    tanh    asin    acos    atan    atan2   sqrt    sin cos tan ceil    floor   fabs    modf    ldexp   _cabs   _hypot  fmod    frexp   _y0 _y1 _yn _logb   _nextafter          ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n B y t e s ) )   >   0                         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ t c s c p y _ s . i n l                   s t r c p y _ s         ( ( ( _ S r c ) ) )   ! =   N U L L             B u f f e r   i s   t o o   s m a l l           ( L " B u f f e r   i s   t o o   s m a l l "   & &   0 )               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f i l e n o . c                   _ f i l e n o           ( f h   > =   0   & &   ( u n s i g n e d ) f h   <   ( u n s i g n e d ) _ n h a n d l e )                     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ c l o s e . c                     _ c l o s e     ( _ o s f i l e ( f h )   &   F O P E N )               ( " I n v a l i d   f i l e   d e s c r i p t o r .   F i l e   p o s s i b l y   c l o s e d   b y   a   d i f f e r e n t   t h r e a d " , 0 )                                   s t r e a m   ! =   N U L L         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ f r e e b u f . c                       ( f i l e d e s   > =   0   & &   ( u n s i g n e d ) f i l e d e s   <   ( u n s i g n e d ) _ n h a n d l e )                         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ c o m m i t . c                   _ c o m m i t       ( _ o s f i l e ( f i l e d e s )   &   F O P E N )                 f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ w r i t e . c                     _ w r i t e     ( b u f   ! =   N U L L )           _ w r i t e _ n o l o c k           ( ( c n t   &   1 )   = =   0 )         i s l e a d b y t e ( _ d b c s B u f f e r ( f h ) )                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ f i l b u f . c                     _ f i l b u f       f:\dd\vctools\crt\crtw32\lowio\ioinit.c         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f t e l l i 6 4 . c                   _ f t e l l i 6 4           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ f l s b u f . c                         ( " i n c o n s i s t e n t   I O B   f i e l d s " ,   s t r e a m - > _ p t r   -   s t r e a m - > _ b a s e   > =   0 )                             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ l s e e k i 6 4 . c                   _ l s e e k i 6 4           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ g e t b u f . c                     f:\dd\vctools\crt\crtw32\stdio\_getbuf.c            ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n W o r d s ) )   >   0                     w c s c p y _ s             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ s w p r i n t f . c                   _ s w p r i n t f       f:\dd\vctools\crt\crtw32\misc\winsig.c          ( " I n v a l i d   s i g n a l   o r   e r r o r " ,   0 )                 f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ w i n s i g . c                     s i g n a l     r a i s e       U S E R 3 2 . D L L         MessageBoxW     GetActiveWindow     GetLastActivePopup      GetUserObjectInformationW       GetProcessWindowStation         n R p t T y p e   > =   0   & &   n R p t T y p e   <   _ C R T _ E R R C N T                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ d b g r p t t . c                   _ C r t S e t R e p o r t M o d e               f M o d e   = =   _ C R T D B G _ R E P O R T _ M O D E   | |   ( f M o d e   &   ~ ( _ C R T D B G _ M O D E _ F I L E   |   _ C R T D B G _ M O D E _ D E B U G   |   _ C R T D B G _ M O D E _ W N D W ) )   = =   0                                                 _ C r t S e t R e p o r t F i l e           _ V C r t D b g R e p o r t A               _ i t o a _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   Second Chance Assertion Failed: File            <file unknown>      , Line      s t r c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                   _CrtDbgReport: String too long or IO Error              s t r c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   " A s s e r t i o n   f a i l e d :   "   :   " A s s e r t i o n   f a i l e d ! " )                                     Assertion failed:       Assertion failed!           s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ r " )                          s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ n " )                   %s(%d) : %s     s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                     s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                           e   =   m b s t o w c s _ s ( & r e t ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               w c s c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                         _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g                             _ V C r t D b g R e p o r t W           _ i t o w _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )                   S e c o n d   C h a n c e   A s s e r t i o n   F a i l e d :   F i l e                     < f i l e   u n k n o w n >         ,   L i n e         
   w c s c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )                                 w c s c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   L " A s s e r t i o n   f a i l e d :   "   :   L " A s s e r t i o n   f a i l e d ! " )                                     A s s e r t i o n   f a i l e d :               A s s e r t i o n   f a i l e d !               w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )                         w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ r " )                        w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ n " )                 % s ( % d )   :   % s           w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )                           w c s t o m b s _ s ( ( ( v o i d   * ) 0 ) ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                                 s t r c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )                                           _CrtDbgReport: String too long or Invalid characters in String                  w c s t o m b s _ s ( & r e t ,   s z a O u t M e s s a g e ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )                               ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . l o c a l e   ! =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . r e f c o u n t   ! =   N U L L ) )   | |   ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . l o c a l e   = =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . r e f c o u n t   = =   N U L L ) )                                                                                         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ l o c a l r e f . c                     ���    f:\dd\vctools\crt\crtw32\mbstring\mbctype.c         c   > =   - 1   & &   c   < =   2 5 5               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ i s c t y p e . c                     p B l o c k   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h e a p \ e x p a n d . c                     _ e x p a n d _ b a s e         0�D�T�    ... _ C r t S e t R e p o r t H o o k 2             _ _ c r t M e s s a g e W i n d o w A               s t r c p y _ s ( s z E x e N a m e ,   2 6 0 ,   " < p r o g r a m   n a m e   u n k n o w n > " )                         <program name unknown>      D e b u g   % s ! 
 
 P r o g r a m :   % h s % s % s % h s % s % h s % s % h s % s % s % h s % s 
 
 ( P r e s s   R e t r y   t o   d e b u g   t h e   a p p l i c a t i o n ) 
                                         f:\dd\vctools\crt\crtw32\startup\tidtable.c         p n h   = =   0         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h e a p \ h a n d l e r . c p p                   Sun Mon Tue Wed Thu Fri Sat Sunday  Monday  Tuesday     Wednesday   Thursday    Friday  Saturday    Jan Feb Mar Apr May Jun Jul Aug Sep Oct Nov Dec January     February    March   April   June    July    August  September   October     November    December    AM  PM  MM/dd/yy    dddd, MMMM dd, yyyy     HH:mm:ss    S u n       M o n       T u e       W e d       T h u       F r i       S a t       S u n d a y     M o n d a y     T u e s d a y       W e d n e s d a y       T h u r s d a y         F r i d a y     S a t u r d a y         J a n       F e b       M a r       A p r       M a y       J u n       J u l       A u g       S e p       O c t       N o v       D e c       J a n u a r y       F e b r u a r y         M a r c h       A p r i l       J u n e     J u l y     A u g u s t     S e p t e m b e r       O c t o b e r       N o v e m b e r         D e c e m b e r         A M     P M     M M / d d / y y         d d d d ,   M M M M   d d ,   y y y y           H H : m m : s s         _ c r t h e a p         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h e a p \ h e a p i n i t . c                     p N o d e - > _ N e x t   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ e h \ t y p n a m e . c p p                   t y p e _ i n f o : : _ N a m e _ b a s e               s t r c p y _ s   ( ( c h a r   * ) ( ( t y p e _ i n f o   * ) _ T h i s ) - > _ M _ d a t a ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                                 t y p e _ i n f o : : _ N a m e _ b a s e _ i n t e r n a l                     s t r c p y _ s   ( p T m p T y p e N a m e ,   l e n + 2 ,   ( c h a r   * ) p T m p U n d N a m e )                       b u f   ! =   N U L L       f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ c o n v \ c v t . c                 _ c f t o e 2 _ l       s i z e I n B y t e s   >   0               s i z e I n B y t e s   >   ( s i z e _ t ) ( 3   +   ( n d e c   >   0   ?   n d e c   :   0 )   +   5   +   1 )                               s t r c p y _ s ( p ,   ( s i z e I n B y t e s   = =   ( s i z e _ t ) - 1   ?   s i z e I n B y t e s   :   s i z e I n B y t e s   -   ( p   -   b u f ) ) ,   " e + 0 0 0 " )                                       e+000   _ c f t o e _ l         _ c f t o a _ l         s i z e I n B y t e s   >   ( s i z e _ t ) ( 1   +   4   +   n d e c   +   6 )                     _ c f t o f 2 _ l       _ c f t o f _ l         _ c f t o g _ l             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t a r t u p \ i 3 8 6 \ f p 8 . c                       _ s e t d e f a u l t p r e c i s i o n             _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   0 x 0 0 0 1 0 0 0 0 ,   0 x 0 0 0 3 0 0 0 0 )                         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          �      	                                   f:\dd\vctools\crt\crtw32\startup\stdargv.c          f:\dd\vctools\crt\crtw32\startup\stdenvp.c          f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t a r t u p \ s t d e n v p . c                     _ s e t e n v p         s t r c p y _ s ( * e n v ,   c c h a r s ,   p )               f:\dd\vctools\crt\crtw32\misc\a_env.c           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ v s p r i n t f . c                   _ v s n p r i n t f _ l             ( c o u n t   = =   0 )   | |   ( s t r i n g   ! =   N U L L )                        ���5�h!����?      �?                            �?5�h!���>@�������             ��      �@      �                            �}    �H�}���E�}���M�}���-�}���\~��g'                L C _ A L L     L C _ C O L L A T E         L C _ C T Y P E         L C _ M O N E T A R Y       L C _ N U M E R I C         L C _ T I M E       	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~                         ( " I n v a l i d   p a r a m e t e r   f o r   _ c o n f i g t h r e a d l o c a l e " , 0 )                           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ w s e t l o c a . c                     _ c o n f i g t h r e a d l o c a l e           f:\dd\vctools\crt\crtw32\misc\wsetloca.c            L C _ M I N   < =   _ c a t e g o r y   & &   _ c a t e g o r y   < =   L C _ M A X                     _ w s e t l o c a l e       = ;     ;   _ w s e t l o c a l e _ n o l o c k             w c s n c p y _ s ( l c t e m p ,   ( s i z e o f ( l c t e m p )   /   s i z e o f ( l c t e m p [ 0 ] ) ) ,   s ,   l e n )                               _ w s e t l o c a l e _ s e t _ c a t               w c s c p y _ s ( p c h _ c a t _ l o c a l e ,   c c h ,   l c t e m p )                   =   _ w s e t l o c a l e _ g e t _ a l l           w c s c a t _ s ( p c h ,   c c h ,   L " ; " )             _ e x p a n d l o c a l e           w c s n c p y _ s ( l o c a l e N a m e O u t p u t ,   l o c a l e N a m e S i z e I n C h a r s , _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   ( s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   /   s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e [ 0 ] ) ) )                                                                             w c s c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   L " C " )                   C       w c s n c p y _ s ( l o c a l e N a m e O u t p u t ,   l o c a l e N a m e S i z e I n C h a r s ,   n a m e s . s z L o c a l e N a m e ,   w c s l e n ( n a m e s . s z L o c a l e N a m e )   +   1 )                                             w c s n c p y _ s ( c a c h e o u t ,   c a c h e o u t L e n ,   e x p r ,   c h a r a c t e r s I n E x p r e s s i o n   +   1 )                             w c s n c p y _ s ( l o c a l e N a m e O u t p u t ,   l o c a l e N a m e S i z e I n C h a r s ,   e x p r ,   c h a r a c t e r s I n E x p r e s s i o n   +   1 )                                         w c s n c p y _ s ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   ( s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   /   s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e [ 0 ] ) ) ,   e x p r ,   c h a r a c t e r s I n E x p r e s s i o n   +   1 )                                                                         w c s n c p y _ s ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   ( s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   /   s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e [ 0 ] ) ) ,   l o c a l e N a m e O u t p u t ,   w c s l e n ( l o c a l e N a m e O u t p u t )   +   1 )                                                                             w c s n c p y _ s ( c a c h e i n ,   c a c h e i n L e n ,   e x p r ,   c h a r a c t e r s I n E x p r e s s i o n   +   1 )                                 w c s c p y _ s ( o u t p u t ,   s i z e I n C h a r s ,   c a c h e o u t )                   _ w c s c a t s         w c s c a t _ s ( o u t s t r ,   n u m b e r O f E l e m e n t s ,   (   * ( w c h a r _ t   *   * ) ( ( s u b s t r   + =   (   ( s i z e o f ( w c h a r _ t   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   -   (   ( s i z e o f ( w c h a r _ t   * )   +   s i z e o f ( i n t )   -   1 )   &   ~ ( s i z e o f ( i n t )   -   1 )   ) )   ) )                                                                                   _ _ l c _ w c s t o l c         w c s n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   & w l o c a l e [ 1 ] ,   1 6 - 1 )                                               _ . ,       w c s n c p y _ s ( n a m e s - > s z L a n g u a g e ,   ( s i z e o f ( n a m e s - > s z L a n g u a g e )   /   s i z e o f ( n a m e s - > s z L a n g u a g e [ 0 ] ) ) ,   w l o c a l e ,   l e n )                                             w c s n c p y _ s ( n a m e s - > s z C o u n t r y ,   ( s i z e o f ( n a m e s - > s z C o u n t r y )   /   s i z e o f ( n a m e s - > s z C o u n t r y [ 0 ] ) ) ,   w l o c a l e ,   l e n )                                           w c s n c p y _ s ( n a m e s - > s z C o d e P a g e ,   ( s i z e o f ( n a m e s - > s z C o d e P a g e )   /   s i z e o f ( n a m e s - > s z C o d e P a g e [ 0 ] ) ) ,   w l o c a l e ,   l e n )                                             _ _ l c _ l c t o w c s         w c s c p y _ s ( l o c a l e ,   n u m b e r O f E l e m e n t s ,   n a m e s - > s z L a n g u a g e )                           _   .   _ _ c o p y _ l o c a l e _ n a m e                 w c s n c p y _ s ( l o c a l e N a m e C o p y ,   c c h + 1 ,   l o c a l e N a m e ,   c c h + 1 )                       s   ! =   N U L L           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ m b s t o w c s . c                       _ m b s t o w c s _ l _ h e l p e r                 ( p w c s   = =   N U L L   & &   s i z e I n W o r d s   = =   0 )   | |   ( p w c s   ! =   N U L L   & &   s i z e I n W o r d s   >   0 )                               _ m b s t o w c s _ s _ l           b u f f e r S i z e   < =   I N T _ M A X           r e t s i z e   < =   s i z e I n W o r d s             p w c s   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ w c s t o m b s . c                       _ w c s t o m b s _ l _ h e l p e r                 ( d s t   ! =   N U L L   & &   s i z e I n B y t e s   >   0 )   | |   ( d s t   = =   N U L L   & &   s i z e I n B y t e s   = =   0 )                               _ w c s t o m b s _ s _ l           s i z e I n B y t e s   >   r e t s i z e           f:\dd\vctools\crt\crtw32\stdio\stream.c         ccs UTF-8   UTF-16LE    UNICODE         f i l e n a m e   ! =   N U L L         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ o p e n . c                     m o d e   ! =   N U L L         ( " I n v a l i d   f i l e   o p e n   m o d e " , 0 )                 _ o p e n f i l e       ( * m o d e   = =   _ T ( ' \ 0 ' ) )           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f t e l l . c                     f t e l l       _ f t e l l _ n o l o c k               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ l s e e k . c                     _ l s e e k     ( " I n v a l i d   f i l e   d e s c r i p t o r " , 0 )               c c s   U T F - 8   U T F - 1 6 L E     U N I C O D E               _ w o p e n f i l e         _ v s p r i n t f _ l       _ v s c p r i n t f _ h e l p e r           _ v s n p r i n t f _ h e l p e r           f o r m a t   ! =   N U L L         _ v s p r i n t f _ s _ l               s t r i n g   ! =   N U L L   & &   s i z e I n B y t e s   >   0                   ( " B u f f e r   t o o   s m a l l " ,   0 )               _ v s n p r i n t f _ s _ l         (null)  ( n u l l )                EEE50 P    ( 8PX 700WP        `h````  xpxxxx                              f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ o u t p u t . c                   _ o u t p u t _ l       ( c h   ! =   _ T ( ' \ 0 ' ) )         ( " ' n '   f o r m a t   s p e c i f i e r   d i s a b l e d " ,   0 )                 f:\dd\vctools\crt\crtw32\stdio\output.c         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ w c s i c m p . c                   _ w c s i c m p _ l         _ w c s i c m p         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ t i m e \ t z s e t . c                   _ t z s e t _ n o l o c k           _ g e t _ t i m e z o n e ( & t i m e z o n e )             _ g e t _ d a y l i g h t ( & d a y l i g h t )             _ g e t _ d s t b i a s ( & d s t b i a s )             TZ  f:\dd\vctools\crt\crtw32\time\tzset.c               s t r c p y _ s ( l a s t T Z ,   s t r l e n ( T Z )   +   1 ,   T Z )                 s t r n c p y _ s ( t z n a m e [ 0 ] ,   6 4 ,   T Z ,   3 )                   s t r n c p y _ s ( t z n a m e [ 1 ] ,   6 4 ,   T Z ,   3 )               c v t d a t e       _ i s i n d s t _ n o l o c k           SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec                ( _ D a y l i g h t   ! =   N U L L )               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ t i m e \ t i m e s e t . c                   _ g e t _ d a y l i g h t               ( _ D a y l i g h t _ s a v i n g s _ b i a s   ! =   N U L L )                 _ g e t _ d s t b i a s         ( _ T i m e z o n e   ! =   N U L L )           _ g e t _ t i m e z o n e               ( _ B u f f e r   ! =   N U L L   & &   _ S i z e I n B y t e s   >   0 )   | |   ( _ B u f f e r   = =   N U L L   & &   _ S i z e I n B y t e s   = =   0 )                                   _ g e t _ t z n a m e       _ R e t u r n V a l u e   ! =   N U L L             _ I n d e x   = =   0   | |   _ I n d e x   = =   1             M S V C R 1 2 0 D . d l l   b i n \ M S P D B 1 2 0 . D L L                          ���   ��� �  A D V A P I 3 2 . D L L         RegOpenKeyExW   RegQueryValueExW    RegCloseKey         S O F T W A R E \ M i c r o s o f t \ V i s u a l S t u d i o \ 1 2 . 0 \ S e t u p \ V C                       P r o d u c t D i r         D L L       M S P D B 1 2 0         M S P D B 1 2 0         PDBOpenValidate5        f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ t c s c a t _ s . i n l                   w c s c a t _ s         S t r i n g   i s   n o t   n u l l   t e r m i n a t e d               ( L " S t r i n g   i s   n o t   n u l l   t e r m i n a t e d "   & &   0 )                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ t c s n c p y _ s . i n l                     w c s n c p y _ s       ( " I n v a l i d   e r r o r _ m o d e " ,   0 )                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ e r r m o d e . c                   _ s e t _ e r r o r _ m o d e           s t r n c p y _ s       _ R a n d o m V a l u e   ! =   N U L L                 f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ r a n d _ s . c                     r a n d _ s     ( " r a n d _ s   i s   n o t   a v a i l a b l e   o n   t h i s   p l a t f o r m " ,   0 )                       SystemFunction036           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ _ s f t b u f . c                     f:\dd\vctools\crt\crtw32\stdio\_sftbuf.c            f l a g   = =   0   | |   f l a g   = =   1             f:\dd\vctools\crt\crtw32\lowio\osfinfo.c                f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ o s f i n f o . c                     _ g e t _ o s f h a n d l e         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ i s a t t y . c                   _ i s a t t y           _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   1   | |   _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   2                                                 f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ m b t o w c . c                       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ r e a d . c                   _ r e a d       ( c n t   < =   I N T _ M A X )         _ r e a d _ n o l o c k         ( i n p u t b u f   ! =   N U L L )             f:\dd\vctools\crt\crtw32\lowio\read.c               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ v s w p r i n t . c                   _ v s w p r i n t f _ l         _ v s c w p r i n t f _ h e l p e r             _ v s w p r i n t f _ h e l p e r           _ v s w p r i n t f _ s _ l             s t r i n g   ! =   N U L L   & &   s i z e I n W o r d s   >   0                   _ v s n w p r i n t f _ s _ l           _ w o u t p u t _ l         s t r c a t _ s         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ x t o a . c                   x t o a _ s     s i z e I n T C h a r s   >   0         s i z e I n T C h a r s   >   ( s i z e _ t ) ( i s _ n e g   ?   2   :   1 )                   2   < =   r a d i x   & &   r a d i x   < =   3 6               l e n g t h   <   s i z e I n T C h a r s           x 6 4 t o a _ s         x t o w _ s     x 6 4 t o w _ s         f:\dd\vctools\crt\crtw32\misc\initmon.c         p l o c i - > l c o n v _ m o n _ r e f c o u n t   >   0                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ i n i t m o n . c                   f:\dd\vctools\crt\crtw32\misc\initnum.c         p l o c i - > l c o n v _ n u m _ r e f c o u n t   >   0               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ i n i t n u m . c                   f:\dd\vctools\crt\crtw32\misc\inittime.c                p l o c i - > l c _ t i m e _ c u r r - > r e f c o u n t   >   0                       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ i n i t t i m e . c                         ��ȴԴ������(�0�<�L�\��Qh�p�|�����������������4p����������������ĵȵ̵еԵصܵ����������� �������$�0�<�H�d�p�����ж���<�h�����ط�(�<�@�H�\���������и��$�P�����Թ��(�\����Q��̺��,�                                                                                __based(    __cdecl     __pascal    __stdcall   __thiscall      __fastcall      __vectorcall    __clrcall   __eabi  __ptr64     __restrict      __unaligned     restrict(    new     delete     =   >>  <<  !   ==  !=  []  operator    ->  ++  --  +   &   ->* /   %   <   <=  >   >=  ,   ()  ~   ^   |   &&  ||  *=  +=  -=  /=  %=  >>= <<= &=  |=  ^=  `vftable'   `vbtable'   `vcall'     `typeof'    `local static guard'        `string'    `vbase destructor'      `vector deleting destructor'        `default constructor closure'       `scalar deleting destructor'        `vector constructor iterator'       `vector destructor iterator'        `vector vbase constructor iterator'         `virtual displacement map'      `eh vector constructor iterator'        `eh vector destructor iterator'         `eh vector vbase constructor iterator'          `copy constructor closure'      `udt returning'     `EH `RTTI   `local vftable'     `local vftable constructor closure'          new[]   delete[]   `omni callsig'      `placement delete closure'      `placement delete[] closure'        `managed vector constructor iterator'           `managed vector destructor iterator'        `eh vector copy constructor iterator'           `eh vector vbase copy constructor iterator'         `dynamic initializer for '      `dynamic atexit destructor for '        `vector copy constructor iterator'          `vector vbase copy constructor iterator'            `managed vector copy constructor iterator'          `local static thread guard'          Type Descriptor'        Base Class Descriptor at (          Base Class Array'       Class Hierarchy Descriptor'         Complete Object Locator'       CV:     ::  template-parameter-     generic-type-   `   '   `anonymous namespace'       ''  `non-type-template-parameter        void    `template-parameter     NULL    }'  }'  `vtordispex{    `vtordisp{      `adjustor{      `local static destructor helper'        `template static data member constructor helper'            `template static data member destructor helper'             static      virtual     private:    protected:      public:     [thunk]:    extern "C"      )   char    short   int     long    unsigned    void    volatile    std::nullptr_t      <ellipsis>      ,...    ,<ellipsis>      throw(     cpu amp ,   char    short   int long    float   double  bool    __int8  __int16     __int32     __int64     __int128    <unknown>   wchar_t     __w64   UNKNOWN     signed      const    volatile   `unknown ecsu'      union   struct      class   coclass     cointerface     enum    volatile    const   cli::array<     cli::pin_ptr<   )[  {flat}  {for    s   .�_�_�_    d.�j�m6    �.�kLB�?    /�Y�>�j    x/B[�M\s    �/�\�N�=     ??     f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ _ f p t o s t r . c                       _ f p t o s t r             s i z e I n B y t e s   >   ( s i z e _ t ) ( ( d i g i t s   >   0   ?   d i g i t s   :   0 )   +   1 )                           p f l t   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ c o n v \ c f o u t . c                 _ f l t o u t 2         s t r c p y _ s ( r e s u l t s t r ,   r e s u l t s i z e ,   a u t o f o s . m a n )                         ( o p t i o n s   &   ~ _ T W O _ D I G I T _ E X P O N E N T )   = =   0                       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ o u t p u t f o r m a t . c                       _ s e t _ o u t p u t _ f o r m a t             ( " I n v a l i d   i n p u t   v a l u e " ,   0 )             f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ t r a n \ c o n t r l f p . c                   _ c o n t r o l f p _ s         �E N U   (�E N U   P�E N U   x�E N A   ��N L B   ��E N C   ��Z H H   ��Z H I   ��C H S   ��Z H H   �C H S   D�Z H I   p�C H T   ��N L B   ��E N U   ��E N A   �E N L   ,�E N C   H�E N B   t�E N I   ��E N J   ��E N Z   ��E N S   �E N T   H�E N G   d�E N U   ��E N U   ��F R B   ��F R C   ��F R L   �F R S   4�D E A   \�D E C   ��D E L   ��D E S   ��E N I   ��I T S    �N O R   8�N O R   `�N O N   ��P T B   ��E S S   ��E S B   �E S L   8�E S O   `�E S C   ��E S D   ��E S F   ��E S E   (�E S G   T�E S H   |�E S M   ��E S N   ��E S I   ��E S A   �E S Z   @�E S R   `�E S U   ��E S Y   ��E S V   ��S V F   �D E S   �E N G   �E N U   $�E N U                                                                                                                                                               a m e r i c a n         a m e r i c a n   e n g l i s h         a m e r i c a n - e n g l i s h         a u s t r a l i a n         b e l g i a n       c a n a d i a n         c h h       c h i       c h i n e s e       c h i n e s e - h o n g k o n g         c h i n e s e - s i m p l i f i e d             c h i n e s e - s i n g a p o r e           c h i n e s e - t r a d i t i o n a l           d u t c h - b e l g i a n           e n g l i s h - a m e r i c a n         e n g l i s h - a u s       e n g l i s h - b e l i z e         e n g l i s h - c a n       e n g l i s h - c a r i b b e a n           e n g l i s h - i r e       e n g l i s h - j a m a i c a           e n g l i s h - n z         e n g l i s h - s o u t h   a f r i c a             e n g l i s h - t r i n i d a d   y   t o b a g o               e n g l i s h - u k         e n g l i s h - u s         e n g l i s h - u s a       f r e n c h - b e l g i a n         f r e n c h - c a n a d i a n           f r e n c h - l u x e m b o u r g           f r e n c h - s w i s s         g e r m a n - a u s t r i a n           g e r m a n - l i c h t e n s t e i n           g e r m a n - l u x e m b o u r g           g e r m a n - s w i s s         i r i s h - e n g l i s h           i t a l i a n - s w i s s           n o r w e g i a n       n o r w e g i a n - b o k m a l         n o r w e g i a n - n y n o r s k           p o r t u g u e s e - b r a z i l i a n             s p a n i s h - a r g e n t i n a           s p a n i s h - b o l i v i a           s p a n i s h - c h i l e           s p a n i s h - c o l o m b i a         s p a n i s h - c o s t a   r i c a             s p a n i s h - d o m i n i c a n   r e p u b l i c             s p a n i s h - e c u a d o r           s p a n i s h - e l   s a l v a d o r           s p a n i s h - g u a t e m a l a           s p a n i s h - h o n d u r a s         s p a n i s h - m e x i c a n           s p a n i s h - m o d e r n         s p a n i s h - n i c a r a g u a           s p a n i s h - p a n a m a         s p a n i s h - p a r a g u a y         s p a n i s h - p e r u         s p a n i s h - p u e r t o   r i c o           s p a n i s h - u r u g u a y           s p a n i s h - v e n e z u e l a           s w e d i s h - f i n l a n d           s w i s s       u s     u s a       |�U S A   ��G B R   ��C H N   ��C Z E   ��G B R   ��G B R   ��N L D   �H K G   (�N Z L   D�N Z L   L�C H N   d�C H N   |�P R I   ��S V K   ��Z A F   ��K O R   ��Z A F   �K O R    �T T O   �G B R   L�G B R   p�U S A   �U S A                                                           a m e r i c a       b r i t a i n       c h i n a       c z e c h       e n g l a n d       g r e a t   b r i t a i n           h o l l a n d       h o n g - k o n g       n e w - z e a l a n d       n z     p r   c h i n a         p r - c h i n a         p u e r t o - r i c o       s l o v a k     s o u t h   a f r i c a         s o u t h   k o r e a       s o u t h - a f r i c a         s o u t h - k o r e a       t r i n i d a d   &   t o b a g o           u n i t e d - k i n g d o m         u n i t e d - s t a t e s           A          f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ g e t q l o c . c                   _ _ g e t _ q u a l i f i e d _ l o c a l e             w c s n c p y _ s ( l p O u t S t r - > s z L o c a l e N a m e ,   ( s i z e o f ( l p O u t S t r - > s z L o c a l e N a m e )   /   s i z e o f ( l p O u t S t r - > s z L o c a l e N a m e [ 0 ] ) ) ,   _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   w c s l e n ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   +   1 )                                                                           L a n g C o u n t r y E n u m P r o c E x           w c s n c p y _ s ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   ( s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   /   s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e [ 0 ] ) ) ,   l p L o c a l e S t r i n g ,   w c s l e n ( l p L o c a l e S t r i n g )   +   1 )                                                                         L a n g u a g e E n u m P r o c E x             G e t L o c a l e N a m e F r o m D e f a u l t             w c s n c p y _ s ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e ,   ( s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e )   /   s i z e o f ( _ p s e t l o c _ d a t a - > _ c a c h e L o c a l e N a m e [ 0 ] ) ) ,   l o c a l e N a m e ,   w c s l e n ( l o c a l e N a m e )   +   1 )                                                                     A C P       O C P       6-    ( p a t h   ! =   N U L L )             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ o p e n . c                   _ o p e n       ( p f h   ! =   N U L L )           _ s o p e n _ h e l p e r               ( ( p m o d e   &   ( ~ ( _ S _ I R E A D   |   _ S _ I W R I T E ) ) )   = =   0 )                     s 1   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m b s t r i n g \ m b s n b c m p . c                     _ m b s n b c m p _ l       s 2   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m b s t r i n g \ m b s n b i c m . c                     _ m b s n b i c m p _ l         _ w o p e n     _ w s o p e n _ h e l p e r         CreateFile2     _ w s o p e n _ n o l o c k         _ g e t _ f m o d e ( & f m o d e )             (   " I n v a l i d   o p e n   f l a g "   ,   0   )               (   " I n v a l i d   s h a r i n g   f l a g "   ,   0   )                     ( o f l a g   &   ( _ O _ T E X T   |   _ O _ W T E X T   |   _ O _ U 1 6 T E X T   |   _ O _ U 8 T E X T )   )   ! =   0                           0   & &   " I n t e r n a l   E r r o r "           0   & &   " O n l y   U T F - 1 6   l i t t l e   e n d i a n   &   U T F - 8   i s   s u p p o r t e d   f o r   r e a d s "                               f i r s t   ! =   N U L L           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ w c s n i c m p . c                     _ w c s n i c m p _ l       l a s t   ! =   N U L L         _ w c s n i c m p       _ o u t p u t _ p _ l       ( ( t y p e _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                 ( " I n c o r r e c t   f o r m a t   s p e c i f i e r " ,   0 )                       ( ( w i d t h _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                       _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ w i d t h _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                   ( ( p r e c i s _ p o s   > =   0 )   & &   ( * e n d _ p o s   = =   P O S I T I O N _ C H A R )   & &   ( t y p e _ p o s   <   _ A R G M A X ) )                                     _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ p r e c i s _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                                 ( ( t y p e _ p o s > = 0 )   & &   ( t y p e _ p o s < _ A R G M A X ) )                       _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ s h o r t _ a r g ,   c h ,   f l a g s )                                 _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ p t r _ a r g ,   c h ,   f l a g s )                             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ d o u b l e _ a r g ,   c h ,   f l a g s )                               p a s s   = =   F O R M A T _ O U T P U T _ P A S S             _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ i n t 6 4 _ a r g ,   c h ,   f l a g s )                                 _ t v a l i d a t e _ p a r a m _ r e u s e ( & p o s _ v a l u e [ t y p e _ p o s ] ,   e _ l o n g _ l o n g _ a r g ,   c h ,   f l a g s )                                 ( ( s t a t e   = =   S T _ N O R M A L )   | |   ( s t a t e   = =   S T _ T Y P E ) )                         ( " M i s s i n g   p o s i t i o n   i n   t h e   f o r m a t   s t r i n g " ,   0 )                         ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp                       _ o u t p u t _ s _ l       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ p r i n t f . c                   p r i n t f     s i z e I n B y t e s   < =   I N T _ M A X             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ w c t o m b . c                   _ w c t o m b _ s _ l       ( o p t i o n   ! =   N U L L )         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ g e t e n v . c                     g e t e n v     ( _ t c s n l e n ( o p t i o n ,   _ M A X _ E N V )   <   _ M A X _ E N V )                   _ t c s n l e n ( * s e a r c h   +   l e n g t h   +   1 ,   _ M A X _ E N V )   <   _ M A X _ E N V                       p R e t u r n V a l u e   ! =   N U L L             _ g e t e n v _ s _ h e l p e r         ( b u f f e r   ! =   N U L L   & &   s i z e I n T C h a r s   >   0 )   | |   ( b u f f e r   = =   N U L L   & &   s i z e I n T C h a r s   = =   0 )                                       s t r c p y _ s ( b u f f e r ,   s i z e I n T C h a r s ,   s t r )                   p B u f f e r   ! =   N U L L           _ d u p e n v _ s _ h e l p e r         v a r n a m e   ! =   N U L L           s t r c p y _ s ( * p B u f f e r ,   s i z e ,   s t r )               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ t m a k e p a t h _ s . i n l                     _ w m a k e p a t h _ s         ( ( ( _ P a t h ) ) )   ! =   N U L L           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ h \ t s p l i t p a t h _ s . i n l                       _ w s p l i t p a t h _ s           ( L " I n v a l i d   p a r a m e t e r " ,   0 )               C O N O U T $       _ w o u t p u t _ p _ l         _ w o u t p u t _ s _ l             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ f p u t w c . c                   f p u t w c     _ L o c a l e   ! =   N U L L           f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ i n c l u d e \ s t r g t o l d 1 2 . i n l                     _ _ s t r g t o l d 1 2 _ l             f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ c o n v \ x 1 0 f o u t . c                     $ I 1 0 _ O U T P U T           s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # S N A N " )                 1#SNAN      s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N D " )                   1#IND       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N F " )                   1#INF       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # Q N A N " )                 1#QNAN   f : \ d d \ v c t o o l s \ c r t \ f p w 3 2 \ t r a n \ i 3 8 6 \ i e e e 8 7 . c                     _ s e t _ c o n t r o l f p             _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   n e w c t r l ,   m a s k   &   ~ 0 x 0 0 0 8 0 0 0 0 )                             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ s t r n i c m p . c                     _ s t r n i c m p _ l       c o u n t   < =   I N T _ M A X         _ s t r n i c m p           f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ c h s i z e . c                   _ c h s i z e _ s       ( s i z e   > =   0 )           ( ( m o d e   = =   _ O _ T E X T )   | |   ( m o d e   = =   _ O _ B I N A R Y )   | |   ( m o d e   = =   _ O _ W T E X T )   | |   ( m o d e   = =   _ O _ U 8 T E X T )   | |   ( m o d e   = =   _ O _ U 1 6 T E X T ) )                                                   f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ l o w i o \ s e t m o d e . c                     _ s e t m o d e             ( ( m o d e   = =   _ O _ T E X T )   | |   ( m o d e   = =   _ O _ B I N A R Y )   | |   ( m o d e   = =   _ O _ W T E X T ) )                             _ s e t _ f m o d e         ( p M o d e   ! =   N U L L )           _ g e t _ f m o d e         n p t r   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ s t r t o l . c                   s t r t o x l       i b a s e   = =   0   | |   ( 2   < =   i b a s e   & &   i b a s e   < =   3 6 )                       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t d i o \ v p r i n t f . c                     v p r i n t f _ h e l p e r         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ s t r t o q . c                   s t r t o x q       f:\dd\vctools\crt\crtw32\misc\wtombenv.c                f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m b s t r i n g \ m b s n b i c o . c                     _ m b s n b i c o l l _ l           n   < =   I N T _ M A X         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ w c s t o l . c                   w c s t o x l       f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ w c s t o q . c                   w c s t o x q       f:\dd\vctools\crt\crtw32\convert\wcstoq.c               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ s t r t o d . c                   _ s t r t o d _ l       p o p t i o n   ! =   N U L L               f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m i s c \ s e t e n v . c                     _ _ c r t s e t e n v       e q u a l   -   o p t i o n   <   _ M A X _ E N V                   _ t c s n l e n ( e q u a l   +   1 ,   _ M A X _ E N V )   <   _ M A X _ E N V                     f:\dd\vctools\crt\crtw32\misc\setenv.c              ( " C R T   L o g i c   e r r o r   d u r i n g   s e t e n v " , 0 )                   s t r c p y _ s ( n a m e ,   s t r l e n ( o p t i o n )   +   2 ,   o p t i o n )                     c o p y _ e n v i r o n         s t r c p y _ s ( * n e w e n v p t r ,   e n v p t r S i z e ,   * o l d e n v p t r )                     _ s t r i n g 1   ! =   N U L L             f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ s t r i n g \ s t r n i c o l . c                     _ s t r n i c o l l _ l         _ s t r i n g 2   ! =   N U L L         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ c o n v e r t \ w c s t o d . c                   _ w c s t o d _ l       s t r i n g   ! =   N U L L         f : \ d d \ v c t o o l s \ c r t \ c r t w 3 2 \ m b s t r i n g \ m b s c h r . c                     _ m b s c h r _ l       _ _ w s t r g t o l d 1 2 _ l           H                                                           ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            RSDS6^�5&SdC�§�3��7   C:\Program Files\MAXON\CINEMA 4D R13\plugins\STL_Importer\obj\STL_Importer_Win32_Debug.pdb      ;  ;                                                                                                                                                                                                                                                                                                     H�        ����    @   L                   `    (                ��               �    ��    �       ����    @   �        (�        ����    @   �                   �    �                D�               0    <`    D�       ����    @           d�       ����    @   �                   �    �    d�        ����    @   �                    ���               �     <`    ��       ����    @   �                    Ƚ<               P    X    Ƚ        ����    @   <                  ��               �    ��(    �       ����    @   �        ��              P   �        D�              @           d�              @   �                    X�d               x    �X    X�       ����    @   d            p      ���               �    ���(        ��       ����    @   �                     �,               @    L(     �       ����    @   ,                    ��               �    �    �        ����    @   �        �       ����    @   �                        ��                ��                4�<               P    `��    4�       ����    @   <                    \��               �    ���    \�       ����    @   �                    ���                   $���    ��       ����    @   �                    ��`               t    |    ��        ����    @   `                    ���               �    �L(    ��       ����    @   �                    ��               ,    @�L(    ��       ����    @                       ̿|               �    �|    ̿       ����    @   |                     ��               �    ��|     �       ����    @   �                    4�8               L    \�|    4�       ����    @   8                    l��               �    �@�L(        l�       ����    @   �                    h�                   ,`��    h�       ����    @                       ��h               |    ���    ��       ����    @   h                    (��                ���               �    �    ��        ����    @   �                    ��8               L    T    ��        ����    @   8                    ���               �    �T    ��       ����    @   �                    ��                        �        ����    @   �                    8�D               X    `    8�        ����    @   D                    X��               �    �    X�        ����    @   �                    |��                   T    |�       ����    @   �                    ��P               d    p(    ��       ����    @   P                    ���               �    �(    ��       ����    @   �                    ��                   ,�(    ��       ����    @                       �h               |    ��(    �       ����    @   h                    @��               �    ��(    @�       ����    @   �                    h�(               <    LL(    h�       ����    @   (                    ���               �    �(    ��       ����    @   �                    ���               �    L(    ��       ����    @   �                    ��D               X    h��    ��       ����    @   D                    ��               �    ���    �       ����    @   �                    p�                   (��    p�       ����    @                       ��d               x    ���    ��       ����    @   d                    ���               �    �`��    ��       ����    @   �                    $�(               <    P`��    $�       ����    @   (                    L��               �    ����    L�       ����    @   �                    p��                   ���    p�       ����    @   �                    ��T               h    x��    ��       ����    @   T                     ��               �    ���     �       ����    @   �                    d�               (    8��    d�       ����    @                       ��t               �    ���    ��       ����    @   t                    ���               �    ���    ��       ����    @   �                    ��4                H     X ��    ��       ����    @   4                      ��                �     � ��     �       ����    @   �                     h��                !    !��    h�       ����    @   �                     ��T!               h!    |!���    ��       ����    @   T!                    ���!               �!    �!��    ��       ����    @   �!                     �"               ,"    <"��     �       ����    @   "                    ��x"               �"    �"�"���        ��       ����    @   x"        ��       ����    @   �"                   #    �"���                ��0#               D#    `#�"���        ��       ����    @   0#                    ��#               �#    �#X ��    �       ����    @   �#                    x� $               $    $$��    x�       ����    @    $                    ���"                ��x$               �$    �$��    ��       ����    @   x$                    D��$               �$    �$��    D�       ����    @   �$                    l�8%               L%    \%��    l�       ����    @   8%                    ���%               �%    �%���    ��       ����    @   �%                    ���%               &     &��    ��       ����    @   �%                     �\&               p&    �&��     �       ����    @   \&                    ���&               �&    �&'���        ��       ����    @   �&        ��       ����    @   4'                   H'    '���                ��t'               �'    �''���        ��       ����    @   t'                     ��'               �'    (X ��     �       ����    @   �'                    h�D(               X(    h(��    h�       ����    @   D(                    ��4'                ���(               �(    �(��    ��       ����    @   �(                    ��)               0)    D)���    ��       ����    @   )                    ��)               �)    �)��    �       ����    @   �)                    ���)               �)    *��    ��       ����    @   �)                    ��@*               T*    p*�*���        ��       ����    @   @*        �       ����    @   �*                   �*    �*���                4��*               +    (+�*���        4�       ����    @   �*                    `�d+               x+    �+X ��    `�       ����    @   d+                    ���+               �+    �+��    ��       ����    @   �+                    ��*                H�L                �X,               l,    x,(    �       ����    @   X,                    ,��,               �,    �,(    ,�       ����    @   �,                    P�-               $-    4-�,(    P�       ����    @   -                    |�p-               �-    �-    |�        ����    @   p-                    ���-               �-    �-(    ��       ����    @   �-                    ��$.               8.    @.    ��        ����    @   $.                    ��|.               �.    �.@.    ��       ����    @   |.                    ���.               �.    �.@.    ��       ����    @   �.                    �4/               H/    T/@.    �       ����    @   4/                    4��/               �/    �/@.    4�       ����    @   �/                    X��/                0    0@.    X�       ����    @   �/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �z	            �z	����    ����                  "�   89   |9                            (9              9                            ��	����    ����                  �9"�   �9   �9                                    ��	����    ����                  :"�   $:   4:                                    �	����    ����                  t:"�   �:   �:                                    �	����    ����                  �:"�   �:   �:                                    �	����    ����                  4;"�   D;   T;                                    >�����    ����                  �;"�   �;   �;                                    >�����    ����                  �;"�   <   <                            p(    h<       x<�<         �    ����       9F        H�    ����       �h        �Q    �<       �<=(=x<�<        l�    ����       \7        ��    ����       wI        ��    ����       =        F*    \=       l=�<        �    ����       (C        G$    �=       �=�<       ��    ����       c]        kn    �=       �=>�<        ��    ����       L        ��    ����       zP        &    L>       `>>�<        �    ����       �C        �R    �>       �>>�<        @�    ����       �E        �>    �>       �>x<�<        h�    ����       �D        Jg    $?       4?�<        ��    ����       bh        `    h?       |?x<�<        ��    ����       �;    ����P�"�   �?                           ����`�"�   �?                           �����"�   �?                           ������"�   ,@                           ���� �"�   \@                           ������    ��"�   �@                               ������    ��"�   �@                               ������"�   A                           ������������"�   4A                               "�   �A                       ���������(�����@�����X�����p�        ����P�    X�"�   �A                               ������    ��������"�    B                               ������"�   DB                           "�   �B                       ������������   ��   ��������        ������"�   �B                           �����"�   �B                           ����P�"�   (C                           ������"�   XC                           �����"�   �C                           ����P�"�   �C                           ������"�   �C                           ������    ��"�   D                               ������������   ��   ��"�   TD                               ����@�����K�   S�   ^�"�   �D                               ������"�   �D                           ������    ������"�   E                               ������"�   `E                           ���� ������"�   �E                               ����������   #�   .�"�   �E                               ����@�����H�   P�   X�"�   F                               ���� �"�   dF                           ������"�   �F                           ����`�    {�����{�"�   �F                               @           �u����    ����                  G"�   G   (G                       ����P�"�   hG                           ������"�   �G                           "�   �G                       ��������������������������9�����T�����o������������������������������������                "�   �H                       ���������������#�����>�����Y�����t����������������������������������������1�                �����"�    I                           ���� �"�   0I                           ������    ��������"�   `I                               ������"�   �I                           ����p�    ��������"�   �I                               ������"�   J                           ������    ��������"�   HJ                               ������"�   �J                           ����p�    ��������"�   �J                               ������"�    K                           ������"�   0K                           ����`�"�   `K                           ������"�   �K                           ������"�   �K                           ����p�"�   �K                           ����@�"�    L                           �����"�   PL                           "�
   �L                       �����    �   �   �   �   �   �   �   �   �            @           _H@           �H����    ����                  "�    M   dM                           M               M                ������    ��"�   �M                               ������    ��"�   �M                               ������    ��������"�   N                               ���� �"�   XN                           �����     � "�   �N                               ���� �    ������"�   �N                               ����@�"�   O                           "�   \O                       ������������   ��   ��������        ������"�   �O                           ���� �"�   �O                           ����@�"�   �O                           ������"�   P                           ���� �"�   LP                           ����@�"�   |P                           ������"�   �P                           ����`�    h�"�   �P                               ����`�����k�   s�   ~�"�   Q                               ����@�����K�   S�   ^�"�   dQ                               ���� �"�   �Q                           ������    ��������"�   �Q                               ������"�   $R                           ����  ���� "�   TR                               ���� ������   �   �"�   �R                               ������������   ��   ��"�   �R                               ������"�   (S                           ���� �"�   XS                           ������    ��������"�   �S                               @           D����    ����                  �S"�   �S   �S                       ������"�   ,T                           ����`�"�   \T                           "�   �T                       ������    ��   �������   �        ����@    H   P"�   �T                               ������"�   $U                           ���� �"�   TU                           ������    ��������"�   �U                               ����@�"�   �U                           ������"�   �U                           ������    ��������"�   (V                               �����"�   lV                           ����P�"�   �V                           "�   �V                       ������������������   ��   ��   ��   ��   ��   ��   �   �
   >�   `�   ��   ��   ��   ��   ��   ��   ��                    ������"�   �W                           ������"�   �W                           ����`�    {�����{�"�   X                               ����`�����h�"�   HX                               ����������"�   �X                               "�   �X                       ������    ��    ��    ��   ��   ��   ��   ��   ��   ��   ��   ��   �   �   �                ����`�"�   lY                           ���� �"�   �Y                           ���� �"�   �Y                           @           k�����    ����                  �Y"�   Z   Z                       ���� �    ;�����;�"�   \Z                               ������"�   �Z                           ������    ��������"�   �Z                               ������"�   [                           ����`�"�   D[                           ������    ��������"�   t[                               @           �����    ����                  �["�   �[   �[                       ������"�   \                           ������"�   H\                           ����@�"�   x\                           ���� �"�   �\                           ������"�   �\                           ����@�"�   ]                           ������"�   8]                           ���� �"�   h]                           ������    ��������"�   �]                               �����"�   �]                           "�   0^                       ����P�����[�   c�   n�����v�        ������"�   `^                           ������"�   �^                           �����"�   �^                           ����P�"�   �^                           ������"�    _                           �����"�   P_                           ������"�   �_                           �����    �"�   �_                               ������������   �   �"�   �_                               ������������   ��   ��"�   8`                               ������"�   �`                           ����p�    ��������"�   �`                               ����p�"�   �`                           ������������"�   (a                               ������������   ��   ��"�   da                               ����0�����8�   @�   H�"�   �a                               ����P�"�   �a                           ������"�   ,b                           ����P�    k�����k�"�   \b                               @            ����    ����                  �b"�   �b   �b                       ������"�    c                           ����0�"�   0c                           "�   �c                       ����P�    h�   ������h�   ��        �����     �     "�   �c                               ����P�"�   �c                           ������"�   (d                           ����P�    h�����h�"�   Xd                               �����"�   �d                           ����P�"�   �d                           �����    +�����+�"�   �d                               ������"�   @e                           ������"�   pe                           "�   �e                       ������������������   ��   ��   ��   ��   ��   ��   !�   ,�
   N�   p�   ��   ��   ��   ��   ��   ��   ��                    ����p�"�   xf                           ������"�   �f                           ������    ������"�   �f                               ������������"�   g                               ����p�����x�"�   Xg                               "�   �g                       ������    ��    ��    ��   ��   ��   ��   ��   ��   ��   ��   ��   �   �   �                ����0�"�   @h                           ������"�   ph                           ������"�   �h                           ������"�   �h                           ����P�"�    i                           ���� �"�   0i                           "�
   �i                       �����    �   �   �                &   1            @           /F@           eF����    ����                  "�    j   Dj                           �i              �i                ������    ��"�   |j                               ����0�"�   �j                           ������"�   �j                           ������"�   k                           @           +�����    ����                  Hk"�   Xk   hk                       ����@�    [�����[�"�   �k                               ����`�"�   �k                           ������    ��������"�   l                               ����0�"�   `l                           ����0�"�   �l                           ����0�    K�����K�"�   �l                               @           �����    ����                  m"�   m   $m                       ������"�   dm                           ����P�"�   �m                           �����"�   �m                           ������"�   �m                           ������"�   $n                           �����"�   Tn                           ������    ��"�   �n                               �����    +�����+�"�   �n                               ������"�   o                           ����P     X "�   4o                               ����p�"�   po                           ������"�   �o                           ������"�   �o                           ���� �"�    p                           ����p�"�   0p                           ������"�   `p                           ����P�"�   �p                           ������"�   �p                           ������"�   �p                           �����"�    q                           ������"�   Pq                           �����"�   �q                           ����@�"�   �q                           ������"�   �q                           "�	   4r                       ���� �    �   �   �    �   (�   0�    �   0�            "�	   �r                       ������    ��   ��   ��   ��   ��   ��   ��   ��            ������"�    s                           ����p�"�   0s                           ����@"�   `s                           "�
   �s                       �����    �   �   �   �   �   �   �   �   �            �����    �"�   t                               "�   pt                       ����p����������������������������� ����            ����p"�   �t                           "�   u                       ����0    H   a����H   a        ����0    8   @"�   @u                               �����"�   �u                           �����"�   �u                           �����    ������"�   �u                               �����"�   (v                           �����"�   Xv                           ����     ;����;"�   �v                               ���� "�   �v                           ����@"�   �v                           "�   Pw                       �����
�����
����         !   )   4   ?   a   l
   �   �   �   �   �            ?                    �����"�   x                           ���� "�   4x                           �����    ������"�   dx                               ����������"�   �x                               ����@����H"�   �x                               "�   Dy                       ����                &   .   6   A   L   W   b   m   x   �   �                �����"�   �y                           ���� "�   �y                           ����"�   ,z                           @           [x����    ����                  \z"�   lz   |z                       ����p	    �	�����	"�   �z                               �����"�    {                           ���� 	    	����	"�   0{                               ����P"�   t{                           ����0"�   �{                           �����	    �	�����	"�   �{                               @           �z����    ����                  |"�   (|   8|                       �����"�   x|                           �����"�   �|                           ����"�   �|                           �����"�   }                           �����
"�   8}                           �����"�   h}                           ����`    h"�   �}                               ����P
    k
����k
"�   �}                               ����@"�   ~                           �����    �"�   H~                               �����"�   �~                           ���� "�   �~                           �����"�   �~                           �����"�                              "�	   h                       ����     (   0   8   @   H   P   @   P                ����    ����    ����    0^    ����    ����    ����    t�    ����    ����    ����    ��    ����    ����    ����            ��        ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    >�    ����    ����    ����    k�    ����    ����    ����    ��    ����    ����    ����    1�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    '�    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    3�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    >�    ����    ����    ����    N�    ����    ����    ����    9�    ����    ����    ����    ��    ����    ����    ����!�'�    ����    ����    ����    0�    ����    ����    ����    \    ����    ����    ����s�    ����    ����    ����    }    ����    ����    ����    �?    �?�?        ����    ����    ����    �#    �"�"        ����    ����    ����C3I3    ����    ����    ����e �     @           z%����    ����                  �"�    �   0�                       ����    ����    ����y66        m5    ��       ���<        ��    ����       -H        ����    ����    ����    �c    ����    ����    ����    g    ����    ����    ����    zk    ����    ����    ����    ;o    ����P"�   X�                           ����    ����    ����V�i�    ����    ����    ����(�;�    ����    ����    ����    �    ����    ����    �����0�0    ����    ����    ����    �=    ����    ����    ����    <B    ����    ����    ����    E    ����    d���    ����    �^    ����    ����    ����    �a    ����    ����    ����    q    ����    ����    ����    �t    ����    ����    ����    �    ����    ����    ����    j�    ����    ����    ����    X    ����    ����    ����    v�        ǖ        ����    ���    ����    �        :�        ����    ����    ����    ��    ����    ����    ����    x�    ����    ����    ����    Ѻ    �����"�   �                           ����    ����    ����    ��    ����    ����    ����    �����    r�        ����    ����    ����    M�����    ��        ����    ����    ��������    ����    ����    �����!�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����     -����    9-        ����    ����    ����    _+����    �+        ����    ����    ����    �2        �1        �2            ����    ����    ����    B    ����    ����    ����    �^    ����    ����    ����    =t    ����    ����    ����    �v    ����    ����    ����    T�    ����    ����    ����    5�    ����    ����    ����    ��    ����    ����    ����    H�    ����    ����    �����<�    ����    ����    ����    �        8        ����    ����    ����    ��    ����    ����    ����        ����    ����    ����    �    ����    ����    ����    �    ����    |���    ����    �n    ����    |���    ����    �o    �����"�   H�                           ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    R    ����    ����    ����    \    ����    ����    ����    �c    ����    ����    ����    �d    ����    ����    ����    ��    ����    ����    ����    d&    ����    ����    ����    v+    �����"�   ؍                           ����    ����    ����    �8    ���� "�   (�                           ����P"�   X�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       [ǵZ    ��          �� �� �� aP ��   STL_Importer.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                     �   8   �   �   B     ^  �  �  Q   �   �   �  �  �   D   g   �   -   ����       
       Copyright (c) 1992-2004 by P.J. Plauger, licensed by Dinkumware, Ltd. ALL RIGHTS RESERVED.                                       �              �             �               3              �9               A                                         �              �              �             �              �<              @>              2@                                             �              �             �              �<              @>              2@                                @�    @�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             |���������      ����        N�@���Du�  s�                  sqrt                                                                                                                                                                                                                                                                                                                                                         8�:�    ����   (�.   $�T�T�T�T�T�T�T�T�T�x�X�X�X�X�X�X�X�.                                                        	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                    zU          �      ���������              �           @J   DJ   HJ   LJ   TJ   \J!   dJ   lJ   tJ   |J   �J   �J   �J   �J    �J   �J   �J   �J   �J   �J   �J   �J   �J   �J"   �J#   �J$   �J%   �J&   �J                                                       �D        � 0                �����
                                                                               ����������������                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                                     abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                            X��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                                                                                                                            Pl����   C   �n�n�n�n�n�n�n�n ooo o,o4o@oDoHoLoPoToXo\o`odoholopo|o�o�oPo�o�o�o�o�o�o�o�o�o�o�op       p$p0p<pHpTp`plp|p�p�p�p�p�p�pqqq(q4q@qLqXqdqpq|q�q�q�q�q(q�q�q�q�qr(r@rXr`rhr�r�r`                                                                        8�                                   ��            ��            ��            ��            ��                          (�        8���@���                                                            8�X�    ����            �T�T�T�T�T�T�T�T�T�T        <�            ���    ����        ����            �p     ����    PST                                                             PDT                                                             ���                                �&                                                                                                                                                                                                                                                                       �                            ����   :   Y   w   �   �   �   �     /  M  l  ����   ;   Z   x   �   �   �   �     0  N  m                      ����   ���5      @   �  �   ����                                      �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                                          �                                                                                                                                                                                                                                                                                                                                                        ��    .?AVruntime_error@std@@         ��    .?AVexception@std@@         ��    .?AVfailure@ios_base@std@@          ��    .?AVsystem_error@std@@          ��    .?AV_System_error@std@@         ��    .?AVbad_cast@std@@      ��    .?AVCommandData@@       ��    .?AVBaseData@@      ��    .?AVios_base@std@@      ��    .?AV?$_Iosb@H@std@@         ��    .?AV?$basic_ios@DU?$char_traits@D@std@@@std@@           ��    .?AV?$basic_streambuf@DU?$char_traits@D@std@@@std@@             ��    .?AV?$basic_istream@DU?$char_traits@D@std@@@std@@               ��    .?AV?$basic_filebuf@DU?$char_traits@D@std@@@std@@               ��    .?AV?$basic_ifstream@DU?$char_traits@D@std@@@std@@              ��    .?AV_Facet_base@std@@       ��    .?AVfacet@locale@std@@          ��    .?AVcodecvt_base@std@@          ��    .?AUctype_base@std@@        ��    .?AV?$ctype@D@std@@         ��    .?AVerror_category@std@@        ��    .?AV_Generic_error_category@std@@           ��    .?AV_Iostream_error_category@std@@          ��    .?AV_System_error_category@std@@            ��    .?AV?$codecvt@DDH@std@@         ��    .?AVSimplePlugin@@      ��    .?AVNeighbor@@      ��    .?AVGeSortAndSearch@@       ��    .?AVDisjointNgonMesh@@          ��    .?AVGeToolNode2D@@      ��    .?AVGeToolList2D@@      ��    .?AVGeToolDynArray@@        ��    .?AVGeToolDynArraySort@@        ��    .?AVbad_alloc@std@@         ��    .?AVinvalid_argument@std@@          ��    .?AVlogic_error@std@@       ��    .?AVlength_error@std@@          ��    .?AVout_of_range@std@@          ��    .?AVoverflow_error@std@@        ��    .?AVbad_function_call@std@@         ��    .?AVregex_error@std@@       ��    .?AV_Locimp@locale@std@@        ��    .?AV?$num_get@DV?$istreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                       ��    .?AV?$num_put@DV?$ostreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                   ��    .?AV?$numpunct@D@std@@          ��    .?AV?$codecvt@_WDH@std@@        ��    .?AV?$codecvt@GDH@std@@         ��    .?AV?$ctype@_W@std@@        ��    .?AV?$ctype@G@std@@             ��    .?AV?$num_get@_WV?$istreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                    ��    .?AV?$num_get@GV?$istreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                   ��    .?AV?$numpunct@_W@std@@         ��    .?AUmessages_base@std@@         ��    .?AUmoney_base@std@@        ��    .?AUtime_base@std@@             ��    .?AV?$num_put@_WV?$ostreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                    ��    .?AV?$collate@_W@std@@          ��    .?AV?$messages@_W@std@@         ��    .?AV?$money_get@_WV?$istreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                  ��    .?AV?$money_put@_WV?$ostreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                  ��    .?AV?$moneypunct@_W$0A@@std@@           ��    .?AV?$_Mpunct@_W@std@@          ��    .?AV?$moneypunct@_W$00@std@@            ��    .?AV?$time_get@_WV?$istreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                   ��    .?AV?$time_put@_WV?$ostreambuf_iterator@_WU?$char_traits@_W@std@@@std@@@std@@                   ��    .?AV?$num_put@GV?$ostreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                   ��    .?AV?$numpunct@G@std@@          ��    .?AV?$collate@G@std@@       ��    .?AV?$messages@G@std@@          ��    .?AV?$money_get@GV?$istreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                     ��    .?AV?$money_put@GV?$ostreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                 ��    .?AV?$moneypunct@G$0A@@std@@        ��    .?AV?$_Mpunct@G@std@@       ��    .?AV?$moneypunct@G$00@std@@         ��    .?AV?$time_get@GV?$istreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                      ��    .?AV?$time_put@GV?$ostreambuf_iterator@GU?$char_traits@G@std@@@std@@@std@@                  ��    .?AV?$collate@D@std@@       ��    .?AV?$messages@D@std@@          ��    .?AV?$money_get@DV?$istreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                     ��    .?AV?$money_put@DV?$ostreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                 ��    .?AV?$moneypunct@D$0A@@std@@        ��    .?AV?$_Mpunct@D@std@@       ��    .?AV?$moneypunct@D$00@std@@         ��    .?AV?$time_get@DV?$istreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                      ��    .?AV?$time_put@DV?$ostreambuf_iterator@DU?$char_traits@D@std@@@std@@@std@@                  ��    .?AVbad_typeid@std@@        ��    .?AV__non_rtti_object@std@@         ��    .?AVtype_info@@     ��    .?AVbad_exception@std@@         ��    .?AVDNameNode@@     ��    .?AVcharNode@@      ��    .?AVpcharNode@@     ��    .?AVpDNameNode@@        ��    .?AVDNameStatusNode@@       ��    .?AVpairNode@@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  � � �    0 F \ n � � � � � � �   0 @ L h � � � � � � � 
  & 0 B R f x � � � � � � �   0 B R ^ l ~ � � � � � � �   6 F \ l ~ � � � � � � � � 	 	 4	 J	 d	 ~	 �	 �	 �	 �	 �	 �	 �	 
                                                                                                                 �         (
                        � � �    0 F \ n � � � � � � �   0 @ L h � � � � � � � 
  & 0 B R f x � � � � � � �   0 B R ^ l ~ � � � � � � �   6 F \ l ~ � � � � � � � � 	 	 4	 J	 d	 ~	 �	 �	 �	 �	 �	 �	 �	 
                                                                                                                 %EnterCriticalSection  �LeaveCriticalSection  DeleteCriticalSection !EncodePointer � DecodePointer �WideCharToMultiByte �MultiByteToWideChar �GetStringTypeW  gIsDebuggerPresent mIsProcessorFeaturePresent cGetModuleFileNameW  fGetModuleHandleExW  ;HeapValidate  �GetSystemInfo @RaiseException  �RtlUnwind �GetCommandLineA GetCurrentThreadId  XFatalAppExitA �GetCPInfo �UnhandledExceptionFilter  CSetUnhandledExceptionFilter SetLastError  HInitializeCriticalSectionAndSpinCount � CreateEventW  RSleep 	GetCurrentProcess aTerminateProcess  sTlsAlloc  uTlsGetValue vTlsSetValue tTlsFree �GetStartupInfoW �GetTickCount  gGetModuleHandleW  �GetProcAddress  � CreateSemaphoreW  PGetLastError  GetDateFormatW  �GetTimeFormatW  � CompareStringW  �LCMapStringW  TGetLocaleInfoW  tIsValidLocale �GetUserDefaultLCID  GEnumSystemLocalesW  �LoadLibraryExW  �GetStdHandle  �WriteFile QExitProcess  AreFileApisANSI  CloseHandle �FlushFileBuffers  �GetConsoleCP  �GetConsoleMode  >GetFileType PReadFile  �SetFilePointerEx  �SetConsoleCtrlHandler �OutputDebugStringW  �WaitForSingleObjectEx � CreateThread  �OutputDebugStringA  �WriteConsoleW rIsValidCodePage �GetACP  �GetOEMCP  3HeapFree  6HeapReAlloc 8HeapSize  5HeapQueryInformation  bGetModuleFileNameA  GetCurrentThread  /HeapAlloc �GetProcessHeap  -QueryPerformanceCounter 
GetCurrentProcessId �GetSystemTimeAsFileTime 'GetEnvironmentStringsW  �FreeEnvironmentStringsW �GetTimeZoneInformation  �VirtualQuery  �FreeLibrary "SetStdHandle  NReadConsoleW  � CreateFileW �SetEndOfFile  �SetEnvironmentVariableA KERNEL32.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                                             � 4   �;�;�;�;O<Y<�<=Q=�=�=�>�>!?T?^?�?�?�?�?�?�? � �   060V0v0�0�0�011D1N1v1�1�1�1�1262V2v2�2�2�2$3.3T3^3�3�3�3�34444>4�4�4�4�4�4�4D5N5t5~5�5�5�566D6N6t6~6�6�6�6�6767t7~7�7�7�7�78&8F8f8�8�8�8�89&9F9f9�9�9�9�9:&:F:f:�:�:�:�:;D;N;t;~;�;�;�;�;<6<V<v<�<�<�<�<=6=t=~=�=�=�=�=>&>F>f>s? � D   �34}4�4o56�6:�:�:�:;$;;�;�;�;<<g<�<�<=w=�=�=!>W>�>�> � $   �0�0�0�0i1�2�2�2�2i3�?�?�?�?  	 8   00g0�0�0�0/1C1K1�1�1�1242@2L2�;x<�<�=�=>�>�> 	 4   f0�2364`4�4�6Z7i7y7p8�8�8{9�:�:@;�<�<Q?�?    	 $   P0�0$1�1�23~384�5e6�6�99:�? 0	 4   30�031�1h2�2;4�4�5�5,686�9�9H:�:8;�>?H?T?   @	 D   51?1D1Q1�1�1�12
222272<2Q3x3�3�3�3�3�3V5[5h5u5z5�5�5�5�5   P	 8   2"2i23�3�9�:;0;<;H;T;`;l;x;�;�;�;�;�;�;�;�;�> `	 @   T0�1�2�3�4�4�4�455:5S5g7q7v7�7�7�7�7�7�;�=�=�=�=�=?   p	 H   �0�0[1p1�2h3!4�4�4�4�4a5�5�5�5Q6�6�6�6�9:;;�;�;�;�<#=T=`=�=   �	 (   =0l0x0�0�1:2h2t2�23H3T3�35$6�> �	 8   �1�3 4�5�5$606�7q9�9::�:�:Q;�;<<f<�<=�>�>.? �	    7t7�7t=	>�>�?   �	     _0�0�2Y3�317�:�:�:�:;'; �	     Y3s3)596y7�7�=C>p>|>O?   �	    �2�7*8�8T:�:�:= �	 H   �0�0�0�0�0�0�2�2�2�2�3Q4{4x6�6�6�6�6�6�6�6�677 7�=�=>�>?X?d? �	 ,   �0]1d1�1�1�1t2{2�2{3�3�3�34�4�4�>�?  
 ,   �2�2�2�2�2335�5�5�5�8:@:L:�=�=�? 
 \   0�0�1�1�1�223�3�4�4�4�4�5�5e67�7�7�7�7�8�8u9):L:X:d:;(;�; <<<�<;=�=%>�>-?2?;?�?  
 X   1�1�1P234(444@4L4�4606<6H6T67n8�8�8�8�8o9�9:�:�:P;�;<O<�<L=}=�=f>�>@?q?   0
 \    010�0�0*1/1�1�1	2M2R2�23�34v465�566L7�708�8K9C:h:t:�:G;�;/<�<�<b=�=w>�>�?�?�?   @
 `   m0�0K1�162�2334�45�56}6�6]7�7;8�889�98:�::;�;<�<�<�<�<=�=�=�=>D>J>p>�>�>??�?   P
 T   ?0�091�1B2�2�23 3v3�3Y4�4�56o6�6V7�7M8�8&9�9):�:;};�;?<�<=�=�=f>�>[?�?   `
 h   J0�0&1�1
2z2�2V3�3B4�4"566�6�7�7�7V889\9h9�9W:�:�:�:�:�:6;�;�;<<{<P=t=�=�=!>D>P>\>h>�>M?�?   p
 \   O0�0V1�1O2�273a3�3�3�3�34�45�5�5�6�677o7�7^8�8�9�9�9�:�:�:J;�;B<�<B=�=->�>?�?�? �
 L   o0�0V1�1~2�2Z3�3?4�4*5�56v6�6V7�7c89�9U:�:&;�;�;_<�<r=�=}>�>�?�?   �
 `   "0�0�0�0�01�12�2&3V3�3�3E4l4�4�5�6�6�6w78,8�8�8�89f9s9�9�9�9�9h:�:j;�;=z=�=>�>T?�? �
 X   $0�01z1�12�2�2S3u34{4�45�56&7Y7|7�7�7_8�8%9�9�9O:�:?;�;+<�<={=�=p>?}?�?   �
 H   h0�0h1�1f2�2V3�3F4�4&5Y6|6�6
7v7�7j8�8J9�9-:�:-;�;�;�<9=->�>?�? �
 L   0�01t1�13�3�3�45�5�5d6�6D7�7b89t9�9T:�:4;�;^<�<g=>@>L>�>"?�?   �
 D   R0�0;1�12�2o3�3�3445{5�5[6�78{8�8[9{:�:[;�;?<�<�=k>�>�? �
 T   �0�0�0O1t1�1�12�2�2k3�3K4�4+5�56{6�6Z7�7W8�8K9�9/:�:";�;<�<=�=�=k>�>]?�? �
 <   G0;1�192�2,3�34�4�5�5�677�7K9�9C:�:<�<�<k=�=c>�?   H   !0�0�1f2k2y2383D3�3;4�45�5�5l6�6K7�7,8�89�9�:?;�;T<;=>�>?    D   k0�0k1�1-575A5K5U5_5i5s5}5�5�5�5�5�5�5�5�5�9�9 :�;�;b<=�?     P   b0�0?1�1�1w2�2W3�3K4�4;5�5;6�67�78D9h9t9�9O:�:+;�;<�<=�=�=k>�>?�?   0 P   181D1�1_23�3�3�4�4 5{5�5K6�6+7�78$9H9T9�9B:�:+;<Z<�<�<=t=�>�>�>�?   @ H   $000_1�1�1�2�2�2484D4�4$5�56�6�7�7�7K8�8;9_:�:�:;�;7<�>?{?�? P T   r0�0w1�1k2�2[3�3�4�4�4�4	6,686D6�6�788�89�9:~;�;<D<P<\<'=�=>>�>�>�>�>?�? ` (   0�01�12F3�3?4�4?5�6�6�8/:�:   p @   0�0;2�23{3�4H5�5x6�6?728�8&9�9m:�:�;<z<�<o=�=o>�>�?   � H   .0�0/1�2�2�2?3�5�5�5�5�5
6[6`6w6�9�9�9�9�9�9;�;�;�;�;�;�;�?�?�? � H   00'0q1v1d2i2�3�3�3�344 4P4T4X4\4:9�9(:�:&;�;<�<#=�=->�>?   � D   22�2{3�3�45�5;6�6-7�7"8�89�9�9o:�:�<=�='>�>�>??{?�?   � <   _0�0�12�2K3�3�4k5�5[6�6K7�7�8l:�:�:�:<�<w=+>�>?�? � <   "0�01�1>2�2;3�3�45�5w6�6�78�9R:+<�<=�=>�>?�?   � @   (0�0"1�12�23�344�4
606<6�6/7�7_:�:h;�;�<�<k=�=l>?�? � L   f0�0�1�1{2�2w3�3o4�4h9o9v9}9�9�9�9�9�9�9�9�9�:�<�<�<>0><>�>�>;?�?   �    ;0�0[12�2�8�<        �3    8   �:�:;+;3;9;r;w;�;�;�;�;<<-<5<u<�<�<�<�<�<�<�?   (   0�0�1O2�23o3�3�3�34�788�>�? 0 @   #0�0�12�23�3K4X5�5X6�68�8�9:�:�:o;�;k<�<g=>�>�>_?�? @ \   50K1�182=2o2�233 3�3�3�34�4�4�4D5�576�6F7�7�8�8�8+9�9::+:0:;;;G<�<G=�=O?�?   P L   o0�0o1�1r2�2o3�3o4�4�5O6�677�7J8�8-9�95:�:/;�;<�<={=�=p>�>p?�?   ` H   t0�0_1�1T2�2T3�3K4�4;5�56�67�7�8�9:�:�:w;�;r<=�=>�>?�?�?   p L   �0�0>1�1?2�2�3�3k4�4H5�5+6�67x7�7h8�8h9�9h:�:h;�;h<�<[=�=;>�>?�?�? � P   k0�0K1�1+2�23{3�3[4�4;5�56�6X7|7�7�7b89�9�:�:�:B;�;?<�<?=�=/>�>?�?   � 8   0�01�12{2�2k3�3�4555(545�5B6�6?7�7�8�8�8�8 � ,   �1�1E2J28#838s8�8�8�8�8�899I9Y9m:�: � $   B0`0�344�5�5�5�=�=�=!>&>7> � 4   �1n3�4�4�4�5�5	6�6�6�6\9�9�9�9�9�9�9�=$>0>O? � 8   �1�1�1�1�1�1I2N2a2�3�3�3;4@4S4�9 ::�= >$>(>,>0> �    �071343@3   �    �6H7�788�89�=�=�=        �9�9:�;�;�;�<�?�?    �   C0�0�01Z1�1�1�12M2�2�23@3�3�384\4s4�4�4585h5�5�5�5(6X6�6�6�617l7�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;;; ;$;(;,;0;4;8;<;@;D;�;�;�;#<S<�<�<�<=4=   d   �3�3�3v4�4�4�4�5�5�5�5�68%8@8h8�8�8�8�8S9g9l9t9~9�9F:U:N;�;<%<C<�<�<�<v=�=�=�=�=o>}>d?~?�? 0 X   �0�0�0�0�0�1�13$353�4�4�4=6m6�6�6�6�7�7�7�7�7�7�7�7�7888�9:V;e;�>v?�?�?�?�? @ \   00�0�0�0�061C1]1�12'2/2v2�2�2f3s3�3�34.4�4�4�4<5l5�5�6�687=7�7�78
8F;X;r;�;�;?< P 0   &252p2f3u3�3�4�4�4�5X6v6�6�7�7�8�9<<>   ` $   �0�0g1v1}3W47�8�;�;9<H<�>   p 0   x2�4�45�5�6�6�6&<5<�<�=�=�=�=9>4?�?�?   � H   �0�0�071�1�1�152N2�2�23S3�3�3	4S4l4�8f9u9�9V;e;�;F=U=q=�>�>�>   � @   G0Y0�1�1�2�264E4a46616�7�7�7&989W9=!=�=�=J>R?�?�?�?   � 4   0/0�1�23(3W3v3�4�4g5�5656�6�6�66;E;@=�?   � (   '1�1828b8�8�89B9�9:�:�:d;�>�> � $   �1�1�4�4�7�7�:;g<�<y=�=�>�> � @   3�4�5�5V7e79%96:E:7;Q;<!<�=�=�=�=6>C>]>�>?'?/?v?�?�? � �   60E0g0o0�0�0�0v1�1�1�1�122�2�2�2�263C3]3�34'4/4v4�4�465E5g5o5�5�5�5v6�6�6�6�677�7�7�7�768C8]8�89'9/9v9�9�96:E:g:o:�:�:�:v;�;�;�;�;<<�<�<�<�<6=C=]=�=>'>/>v>�>�>6?E?g?o?�?�?�?   � �   v0�0�0�0�011�1�1�1�162C2]2�23'3/3v3�3�364E4g4o4�4�4�4v5�5�5�5�566�6�6�6�667C7]7�78'8/8v8�8�869E9g9o9�9�9�9v:�:�:�:�:;;�;�;�;�;6<C<]<�<='=/=v=�=�=�>�>?v?�?�?     t   0#0�0�061C1&232�5�5�5F6U6�6�6v7�78%8�89M9�9�9F:U:�:�:v;�;�;<.<�<�<�<=#=N=�=�=�=6>C>n>�>�>�>V?c?�?�?�?    �   0v0�0�011>1�1�1�1&232^2�23S3�3�3�3�3F4S4~4�4�45f5s5�5�56.6�6�6�67#7N7�7�7�768C8n8�8�89�9�9:l:�:L<|<�<�<,=�=�=>L>|>�>�>?<?l?�?�?�?   �   ,0\0�0�0�01L1|12d389=9�9�9�9�9(:-:�:�:�:�:�:�:;	;;�;�;�;�;�;�;<	<<�<�<(=-=�=�=�=>>>->2>7>�>�>�>�>�>??"?'?�?�?�?�? 0 D   11�1�1V2e233�3�3V4e4q5v5�5�5�5�5�5�5�5�6�6�6�6�6�6�6�6�6 @ H   44"4/444@4\4a4f4�4�4�4�4�4 55!5&5f5y5{6�6�7�7�8�8�9G:�?�?�?   P (   .0:0�0�6�6�6777f>u>�>�?�?�?   ` P   �0�001�2�2�2&454p4f5u5�5�6�6�6�7�7-8&959p9f:u:�:�;�;�;�<�<0=&>5>p>f?u?�? p P   �0�0�0�1�102&353p3f4u4�4�5�5�5�6�607&858p8f9u9�9�:�:�:�;�;0<&=5=p=f>u>�> � (   W0�0�0�1�1�2�3�6^8�:�:<<X=9>   �    �0�2F5X5'666�8�9�<? �    F2X2'363�5�6�9<F?U? �     f1u1�3�3+4947&;8;�;�;�> �    �2G5�7�78\9j9�9�9   � (   �0T1�3@7D7H7L7P7�;�;�;L=Z=�=�=   �    �4D5�70;4;8;<;@;�?   � ,   v7�7=8�89�9�9}:0;F;�;W<7=�=�>	?l?     4   &0&191�1V2V3i3�364I4�45%5�5�5�6�676<H<a<    l   �1�1�142M2�2�23a3�3�3!4s4�4�435O5�5�56c6�6�67m7�7�7/8K8�8�89a9�9�9!:q:�:�:1;M;>>Z>�>�>?a?}?�?   \   !0=0�0�0�0S1�1�12c22�2 393�3�3�3M4�4�45a5}5�5!6=6�6�6�6Q7�7�7�:';3;�;�;6=E=�=�=   0 8   �0�0�1�163H3n3�6�6�8�8?? ?$?(?,?�?�?�?�?�?�?   @ 0   63H3n3�6�6�8�8?? ?$?(?,?�?�?�?�?�?�?   P $   �8'9�9�9�9�9�:;�;x<�<�=�>�? ` (   ]0�02,3�3�3|8�8,9C9v<�<�=�=�?�? p <   1%1�2�23�4�4�4�6�6�668E8a8�9�9;;W<i<�=�=�=v?�?�? � 8   1111�2�2�266E6a6&858Q8:%:A:�;�;�;=)=g>y>�?�? � `   1111�2�23f4u4�4�56'6�9�9: :�:M;�<�<=X=�=�>�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   � d    0000022�2�23�3
5G5�5�5467$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8v:�:�:�:   � ,   �122@29�9?:a:�:;;@;&=5=N=p=_?�? � D   0A0�0�0�0 1V2e2~2�2�4*55�57)7�8�8m9�9?:_;�<=�=�=w?�?�?   � @   �1�1�1v4�4�4�4�6�6.7G7Z799s9�9f;u;�;�;�;�=�=7>Q>�>�?   � H   G0c0q0�0�0:2�3�3�3�34w5�5�56�6�6V7h7�7g:�:;!;�;�<=3=A=p=�=
? � P   ^0z0�0�0�0G2X2�2�2w3�3&484U467E7a7w7�7�7�7f9u9�9�9�9�9�9�;<}<�<>�>m?�?   $   �0�0�0v2�2�2�4�4�5�5777�7�7     P1@2�5�5=??        �5�7�7   0 l   24k4G5�5�6�6g8�89%9G9O9�9�9�9V:e:�:�:�:�:�:�;�;�;�;<#<=<�<�<==V=c=}=>%>G>O>�>�>�>V?e?�?�?�?�?�? @ �   �0�0�0�01#1=1�1�122V2c2}2F3S3~3�4�4&535^5�5�5�5F6S6~6�6�67�7�7�7�78v8�8�89L9�9�9�9:L:|:�:=	==#=(=1=J=O=T=>>�>�>V?e?   P `   h0m0z0�0�0�0�0�0�0�3�3444 4<4A4F4�4�4�4&656m6f7u7�7�8�8�8�9�90:&;5;p;f<u<�<�=�=�=�>�> `     1�3�3�35*5�5�5�<=�?   p L   �2�2 333�7�7m8 969V:i:�:6;E;�;�;<d<}<�<=1=�=�=�=6>�>�>�>6?O?�?�? � 0   0V0�0�01c11g3s3�3�3V4b45(5N5�8�8�:�: � D   �0�0 1111l1p1t1x1|1�1�6�6F8U8�9�9v;�;�; <u<-=z>�>�>8?�?   � \   w0�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�3�3404o;�;&<5<N<p<_>�>?%?>?`?   � 0   �0&252�2�2�4�4�4�4
5�6�6�6�6	77�8�89   � (   �0�2�2J6�6�7�8
9z:;)<==T=�>T?   �    y0�1�1(6H6�6};�;�;   �     0�0�0�0)1�1X2�5�67�=   �    3�3�3�3�4�4�4�:�:�?      �7�7:�>  $   <1W1y102�2�34;4�4�488�>        �6�69   0     A0�0E1�2�23�3�3�5a=�=�? @     7�78�9�9�9{:�:?0?L?d? P L    7777O7R<e<�<�<�<�<,=3=@=E=j=�=�=�=�=�=�=�=w>~>�>�>?7?x?}?�?�?�?   ` �   E0J0f0�0�0�0�0�0�0�0�0�0�0�01111#1/181=1C1M1W1i1{1�1�12 2&2,22282?2F2M2T2[2b2i2q2y2�2�2�2�2�2�2�2�2*30363<3B3H3O3V3]3d3k3r3y3�3�3�3�3�3�3�3�3�3!4(4�4�5�6�6�6�6�6�7�7�7�7W9s<�<�<U>s>�>�>�>�>�>�>�>�>?? ?$?(?,?0?4?8?�?�?�?�?�?�? p �   0 0'0,00040U00�0�0�0�0�0�0�0�0�01$1(1,101f4k4t4�4�4�45
55=5B5G5�5�5�5�5�5�5�6�68+898�9::#:+:0:4:8:a:�:�:�:�:�:�:�:�:�:�:;;; ;$;�;�;�;�;�;�;�;�;<A<H<L<P<T<X<\<`<d<�<�<�<�<�<�?   � �   080h0�0�0�0<1|1�12<2l2�25`5e5n5�5�5�5�6�6�6�6�6�6777�9�9�9V:[:m:�:�:�:�:;-;W;k;�;�<�<�<*=/=8=b=g=l=�=�=> >T>Y>b>�>�>�>�?�?�? � �   *0/080b0g0l0�0�01 1T1Y1b1�1�1�1�2�231363;3r3w3�3�3�3�3V4[4m4�4�4�4�4�4�4U5a5�5�5�5�5�5666f7k7}7�7�7�7�7�7�7e8q8�8�8�8�8�89!9&9�:�:�:�:�:�:;; ;J;O;T;�;�;�;*</<8<b<g<l<�<�<�<�<�<�<�=�=�=�?�?�?�?�?�? � �   00"0L0Q0V0�0�0�0�0�0�0Z1_1k1v4{4�4�4�4�4555�5�5�5:6?6H6r6w6|6�6�6�6�6�67Q7V7_7�7�7�7$8A8J8�9�9:#:W:\:e:�:�:�:V<[<m<�<�<�<�<�<�<�=�=�=�=�=�=�=�=�=>>>$>Q>Z>�>�>�>�>??$?T?�?�?�?�? � �   0e0�1�1�1�1�1�122"2Y2^2g2�2�2�2�2P3i3n3z3�3444&4a4j4s4�4�5�5O6_6d6i6n6�6�6�6�6r7~7�7�7�7�7�78)858P8`8l8�8�8�8�8�8C9I9}9�9�9�9�9�9�9�97<H<`<q<f=k=}=�=�=�=/>z>�>�>?1?b?�?�?   � �   <0A061;1M1�133-3H3�3�3�3�3�3�3�34474<4c4�4�4�45N5t5�5�5$6[66�6�6T7X7\7`7�8�8�8�8�8�8999+9H9:;:S:X:�:�:�:�:�:;�;�<�<F=K=]=�=�=�=�=�=�=>>>�>
?.?9? � �   1060B0o0t0y0�0�0�0�0�0�0-121>1k1p1u1
2i3n3z3�3�3�3�3�3 4B4�45%515U5v5{5�5�566�6�6�6�6�6�6
777<7A7N7g7~7�7�7�758A8e8q8�8�89+9\:a:m:�:�:�:�;�;�;<!<&<d<i<u<�<�<�<_=�>�>�>�>4?9?E?r?w?|?�?�?�?�?�? � �   0�0�4&5+5=5z55�5�5�5�5�6�6�667>7G7W7\7h7~7�7�7�7�7�78 8%8U8Z8f8�8�8�8�8�8A9G99�9�9�9:9:?:x:}:�:�:�:�:�:;!;&;L;V;[;g;�;�;�;�;�;�;�;<&>+>=>q>y>�>�>�>�>�>�>�>�>�>�>�>?,?I?N?|?�?�?�?   � �   A0J0�0�0�0�0�0�0�0�0�0�0�0�011S1\1u1�1�263;3M3�3�3�3�3�3�3�3�3�3
44414=4F4l4q4}4�4�4�47�7#8(8-8x8&9+9=9];f;o;;�;�;�;�;�;�;�;�;�;<<9<><x<�<�<==8=X=�=�=�=�=�= >@>N>�>�>�>�>�>�>???#?+?1?:?@?F?M?R?w?�?�?�?�?   �   :0D0I0U0p0�0�0�0�0�0�0�0�0�0�0�2�2B3�4�4�5�5�5�7�7�:�:�<�<=!=/=3=@=D=R=V=d=h=v=z=�=�=�=�=�=�=�=�=>>>f>k>u>�>�>�>�>??d?�?�?�?�?  �   11-1R1u1�122N2c2�3)585G5l5�5�5�566�6�6
77(7d7�7�78>8K8S8[8�8�:`;r;�;�;�;<@<G<t<�<�<�<�<�<=(=5=B=�=�=�=�=�=�=8>[>?(?2?L?�?�?�?�?�?       81h1�1�1�1265F5�599�= 0 $   a0�1f2k2}2�3�3�3l4u4�>�>�>   @     \4j4�4�=>F>�>�>%?e?�?�? P L   %0e0�0Q1V1[1�1�1,2:2�2�2�2�2g3�34*4E4`4�4�7�799"9Y9f9s9�;M<�=�=   ` �   0050A0�0�0�0�0�0�01;1@1E1�1�1�12V2[2`2�233k3�4�45Q5V5_5�5�5�5�5�5�5666E6J6S6}6�6�6�688*8W8\8a8::-:j:o:x:�:�:�:�:�:�:';,;1;I<N<Z<�<�<�<==-=q=v==�=�=�=�=�=�=!>&>+>e>j>s>�>�>�>?   p �  00^0d0�0�0�0�01N1T1�1�1�1�122^2d2�2�2�2�2�23=3C3[3~3�3�3�3�3�34>4D4~4�4�4�4�4�45^5d5t5�5�5�5�56	6E6K6S6]6c6q6v6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67777$7.747B7G7Q7W7e7j7t7z7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 8888#8)878<8F8L8Z8_8i8o8}8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8	9999,919;9A9O9T9^9d9r9w9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9:::!:&:0:6:D:I:S:Y:g:l:v:|:�:�:�:�:�:�:�:�:�:<<6<^<d<�<�<�<�<)=I=i=p=�=�=�=�=�=�=,>Y>T?   � P   '0�0�4�4�45
55F5K5T5~5�5�58*898s8�899*9L9Q9V9�9�9�9�9::u:�:f;u;   � �   +1�1�1�1�1�1�1l3�3�3�3'4,414�5�5�5�5�5�586=6I6v6{6�6�6�6�6
777Z7_7k7�7�7�7�7�78J8T8l8�8�8�:�:�:�:�:+;0;5;�;�;�;�;�;�;V<[<g<�<�<�<===D=I=N=�>�>�>!?&?+?�?�?�?�?�?�? � �   D0I0U0�0�0�0111L1Q1V1�1�1�1�1 22u2z2�2�2�2�2!3&323_3d3i3�344=4B4G4�4�4�4�4�4�4G5L5X5�5�5�5�5�561666;6�6�6�6�6�6�688#8S8X8]8�8�8�8%9*9/9�9�9�9r:w:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;; � \   �1�4�4�4�4�5688 8$8(8,8084888<8@8�8�8�8�8�8�8�8�8;p;u;z;�;�;�;�=�=�=�=P>U>Z>�?   � �   w0|0�0'1,111�1�1�1�2�2�2C3H3M3�3�3�3p4u4z4�455�5�5�5�6�6�6b7g7l7(8-828�8�8�8�9�9�9):.:3:�:�:�:S;X;];R?W?c?�?�?�?�?�?�? � D   0#0(0v0{0�0�0�0�0Z1_1k1�1�1�1�2�2�23
33�7�;$=(=,=0=4=:?   � |   4484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�6D7l7q7}7�8z9�9C:�<�<�=�=>�>�>�>�>f?�?�?�?�?�?�?�? � �   .0400�0�0�01$1m1�1�1�1�12'2N2T2�2�4�45P5�5�5�5"6�6�6�6�6�6�6777<7G7M7S7X7c7�7�7�7�7�7~8�8�8�8�8B9s9�9S:Z:�:,;d;�;�;�;<:<b<�<J=T=�=�=>q>�>�>�>�>�>�>�>?.?8?T?d??�?�?�?   �   E0Q0z0�0A1P1*2J2\2�2�2�2�2�2�2�2�2�2�2X3]3b3i3�3�3�3�3�3�3�3�3�344*5�5�5H6y6~6�6K7�8 9%919^9c9h9�9�9�9�9�9�9
:4:C:Z:�:�:�;�;�;�;�;�;<<<?<D<I<j<�<�<�<�<=�=�=�=�=%>G>N>W>�>�>�>�>�>�>???/?H?M?[?n?�?�?�?�?�?�?�?�?�?�?    �   �0�01!1&1A1N1S1a1i1�1)2.2:2g2l2q2�2�2�2�2�2�2�23�3�3�3�3�3�3�3444K4P4U4m4�4666>6K6W6g6n6�6�6�6�6�6
777 7U7Z7g7l7�7+9�9�9
:+:y:E;?k?     8   M0�0�1�1�2�2�2�23313<3�3�5A6�:~;T<X<\<`<&?h?�? 0 �   060;0M0e0z0�0�102E2Z2�2�2�2�233"3Y4a4�4�4�4�4�455&5<5F5O5?7D7M7w7|7�7�7�788'8Q8V8[8�8�89>9C9L9v9{9�9�9�9�:�:;1;6;;;�;�;�;�;	<<<L<Q<V<|<�<�<�<�<�<�<-=c=h=q=v>�>�>�>?z??�?   @ �   &0+0=0{0�0�0�0�0�0�011161?1i1n1s1�1�1�1222�2�23V3y3~3�3�3�3�3�344%4Z4_4d4�4�4�4�4�5X6]6f6�6�6�6�60757>7v7{7�7�7�7]8g8�859V9m9r9~9�9�9�:�:�;�;�;<`<j<�<=s=�=�>�>?   P `   90C0y0�1�1�1	2'2�2�2�2!3777I7N7S7�8�8�9�9:7:`:�:�:�:1;�;�;�;�;�;�; <�<�<h=�=�=l>x>   ` l   40A0Y0y0�0�0�0�0�0A1F1O1y1~1�1N2_2d2m23�34L4�4�4�5;6D7�8=;B;K;�<�<�<Z=f=�>�>�>0?S?X?a?�?�?�?�?�?�? p �   070<0A0}0�0�0�0�1 2	2;2E2l2�2�2�2�23
33�3�3�3/4=4L4b4�4�4�4�4o5t5}5�5�5�5�5�5M6R6[6�6�6�67!7N7w7|7�7�7�7�7�78�:�:�:;;;L;Q;];�;�;�;D>K>w>�>�>�>�>�>�>�>??#?A?�?�?�? � <  Y0`0g0�0�0�071<1H1u1z11�12*202S2�2�2�2�2�2�2 44V4[4m4�4�4�455A5H5N5U5h5m5t5{5�5�5�5�5�5�5�5�5�5�5>6J6R6s6y6�677D7I7U7�7�7�7�7�7�7�7�7�7�7�8919D9J9Y9g9m9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9::::!:&:,:@:`:g:�:�:�:�:�:�:;;;o;z;�;�;�;�;�;�;4=o=t=�=�=�=�=�=�=�=>>>*>�>�>�>�>�>? ?%?d?i?r?�?�?�?�?�?�?   �   F0K0d0-1K1P1U1}1�1�1�1�1�1�1�1�1J2O2T2�2�2�2�2�2�2�2�2�23#3(3\3m3r3w3|3�3�3�3�34E4J4O4�4�4�4�4�4�4�475<5A5i5n5s5x5�5�5�5M6�67:7I7v7}7�7�7�7�7�7�7}8�:�:�:�;�;�;�;<<2<?<D<J<W<\<b<�<�<�<===#=V=b=n=s=x=�=�=�=�=�=�=>>/>4>9>>>�>�>�>�>????I?N?S?�?�?�?�?�?�?�?   � t   00J0�0T1y1�1�1�1�122)2I2N2S2�2�2
333-373�3�3�34�7m8�9:�:�:�:�<v={=�=�=�=�>?(?b?i?w?�?�?�?�?�?�?�?�? � d   0%0Q0a0k0�0�0�0�1(2z2�2�6�6�6�6757N7W7�8�8�89m9�9�9�9�9:J:|:�:�:�:�:�:�:�;+<�<�<v=�=�=? � �   C0H0Q0�0�0�0�1�1�3�3�3C4J4v4�4�4J5O5X5�5�5�5�5�5�5�56�6�6�7�7�7�7�7�788"8Y8^8g8�8�8�8�8P9i9n9z9�9:::&:a:j:s:�:�;�;M<]<b<g<l<�<�<�<�<m=y=�=�=�=�=�=>$>0>K>[>g>�>�>�>�>�>>?D?x?}?�?�?�?�?�?�?   � �   t1�1�1�1�1�1�2�2A3J3%434G4�4�4�4�45C5�5�5�5�566/7<7B7U7y7�7�7�7848;8Z8_8h8�8�8�8�8�8�8G9`9g9�9�9�9::�:�:�:�:�:;; ;E;�;�;�;�;�;v<{<�<D=J=O=f=k=}=�=�=j>o>t>v?{?�?�? � \   �0�0�0�1�1�1�1�1C2H2Q2�2�23@3J3�3�3�3V4[4m4J5O5�7�7�7�7�7�7*8/8;8h8m8r8�8�8�8999 � �   �1�1�122$2j2o2{2�2�2�233#3P3U3Z3d4i4n4s4h5�677#7P7U7Z7�7�7�7�7�7�7�9�9�9:$:):o:t:�:�:�:�:�<B=G=S=�=�=�=�=�=�=>>>�?�?�?   L   04090>0w0|0�0�0�0�0�6�6�6�6�67�7�7�7�9 :G:_:�:�:�:�:�:�:�:�:$;t;|;  �   X0l0�0�0�0�041X1g1|1�1�1�1�1�1f2q2~2�2�2�2�2�23%33�3�3484[4�4�4�4�4�4�4�5�5�5�5�5�5666D6I6N6�7 8�8<9{:|;�;�;�;�;�;�<�<�<===#=0=�=�=�=>>>�>�>�>(?`?     �   	000q0�0�0�0111f1k1p1�2�2333F3K3P3h3l3p3t34Q4�40555:5�5�5�5�5(6T6Z6777�7�7�7�7�7�7�70858:8v8{8�8�8�8�8H9M9R9�:�:�::;�;F<K<]<�<�=�=K>�>   0 d   70<0A0�0�0�0�0�0151:1?1{12"2g2x2�3.484]4b4g4l4�45h5t596E6�6�6J89�9�9�9%:*:/:�=|>�>�>�>   @ l   �0H12|2�2�2�4 5555 5�586W6�7�7�7�7�7�7�8�8�9�:<<<@<E<J<�<�<=!=-=Z=_=d=�=�=t>{>�>�>�>
???   P �   e0m0�1�1�1�12$2)2`3�3!4�4:6"8'838`8e8j8�8�8,919=9j9o9t9�9�9]:e:�:�:�:�:�:�:�<�<�<�<�< ==Y=q=�=�=�=�=�=>>>N?q?v??�?�?�?�?�?�?   ` �   t0y0�0�0�0�011�2�2�2333J3{3�3�3�3�3�3!4&424_4d4i4�4�4�4I5N5Z5�5�5�5�5�5�56$6)6_6g6�6�6�6�6�6�6�6�6�6�6�6�6�6U9a9l:�:9;>;G;t;y;~;<�<�<1=�=�=�>�>�? p �   +1f3k3}3�3�3�3�3�3�3�4�4�45)5.575l5q5v5�5�5�5�5
666M6�6�6�6�7�7�7�7868@8j8�8�89A9F9O9j9o9x9�9�9�9E:J:S:}:�:�:�:�:�<�<�<�<�<�<=L=Q=]=�=�=�=�=�=>0>5>:>o>�>�>??+?X?]?b?�?�?�?�?�?�?   � X   0080�0�0�0�0�0�0�0�0�0�0�0�0�0z6�6~;�;�;�;+<0<5<�<=@=�=�=�=�=�=�=&>+>4>^>c>h>�? � �   ;0�0�0�01
11L1Q1Z1�1�1�1g3l3x3�3�3�34
44C4H4M4�4�4�4C5�5�566#6P6U6Z6�6�6�7[8�8�8�8999U9Z9f9�9�9�9�9::`:e:q:�:�:�:�:�:
<�<�<�<=	==�=�=�=�=@>E>Q>�>�>�>�>�>�>*?/?4?�? � D   $0S0�0�0�0,1116122[3b3�4�4�5�6C7888B8G8L8T9::J:Q:�:�: � �   �1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1024282<2@2D2H2L2P2T2X2\2`2d2h2�:;;;>;C;H;�;�;�;�;�;�;E=J=S=}=�=�=�=�=�=>
>>   �   00-0B0\0i0q0�0�0�0�1�1�1�1�1�1�1 2222"2*222O2W2_2g2o2{2�2�2�2�2�2�2�2�2�2�2 3333�3�3�3�344)474O4]4�4�4�4666�6�6�6777=7B7G7h7m7r7�7�7�7�7�7�7�7�7�7�788#8-8;8E8U8[8�8�8�89W9_9�9�9�9�9�9�9�9�9 :e:j:o:�;�;�;>>�>�>Q?`?�?�?�?�?�?�?�?�?   � �   000 0&0/070B0L0R0[0d0$141D1T1�1�1�1�1�1�1�1I2N2W2�2�2�2�2	333A3F3K3b3�3�3�3444k4p4y4�4�4�4�4�4�4$5)5.5G5}5�;�;�;�;�;�;<F<h<t<�<:=F=S=a=m=�=�=�=�=�=�=#>D>�>�>�>�>�>�>�> ??1?�? � �   S0m0%1?1�1�1�1�1�1�1�1(2�2�2x33�4�4�4�4�4�455m5r5{5�5�5�5$6,6Y6�6�6�6�6�6�6C7J7w7�7�7�7�7�7�7"8*8�9�9�9�9�9�9;:C:�:�:�: ;	;3;8;=;�;�;�;w<<�<�<�<�<===W=_=�>�>�>�>&?+?4?^?c?h?�?�? � �   00050:0y0�0�0�04191B1l1q1v1�1�1�1�2�2�233393>3C3�3�3�5�5F7K7]7v7G9X9_9�9�9�9�9�9�9�9:::%:S:X:a:�:�:�:�:�:�:�:�:;-;2;7;E;Z;e;p;�;a<f<r<===�=�=�=�=�=)>�>�>�>"?�?�?   �   00-0�0�0�0R1k1�1�1�1�1�12[2s3�3�3�3�3�3�34�4�4�4�4!5&5+5Q5|5�5�5�5�5�5�5f6k6}6�6�6�7�7�7�7�7)8G8#9?9K9t9�9�9�9%:0:i:�:�:�:�:�:�:�:�;�;�;�<=&>+>=>�>�> ??F?K?]?�?�?�?�?  �   000<0g0l0u0�0�0�0�0�0�01161;1t1�1�1�1 3C3H3T3�3�3�3�3�3�3�30454:4t4y4�4�4�4�4�4;5@5L5�5�5�5�5666L6Q6V6�6�6$7)757m7r7w7�7�78>8e8�8�89?9�9�9�9�9:):3::�:�:;];{;�;�;�;<7<=!=+=d=�=l>�>�>?@?v?�?�?   p   =0�0�0�1�1�1�1-2M2k2V3`3j3�3404W4�9M:R:^:�:�:�:@;n;�;=<B<N<{<�<�<�<�<�<�<�<=�>�>?5?:???�?�?�?�?�?�?   0 �   0_0g0�0U1]1�1�1�1�1�1�182?2�34�4�4�4�4�4�4"5'535`5e5j5y7�7P8U8a8�8�8�8�8�8�8999F9�9�9�9�9�9":':,:j:q:�;C<H<T<�<�<�<�<�<�<-=2=7=�=)>X>??   @ t   _0f0�1�1�2�3�4[5`5l5�5�5�5�6a7h7�7�7�7�7 ???????? ?$?(?,?0?4?L?P?T?X?\?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? P �   777G7L7Q7�7�7�7�7�7!8&8+8�8�8�8�8�891969;9�9�9�9:::I:N:S:�:�:<< <M<R<W<�<�<�<�<�<�<==}=�=�=�=�=�=>	>>B>G>L>d?i?u?�?�?�? ` �   �2�2�2333D3I3R3|3�3�3�3�3+40494c4h4m4�4�4�4�4�4�4�5�5�566"6�7�7�7�7�7�70858A8n8s8x8�8�8"9'939`9e9j9�9�9�9�9�9�9;;#;P;U;Z;y>~>�>�>�>�>�>�>?,?1?6?q?y?�?�?�?   p `   00"0a0f0o0�0�0�0�1�1�1�1�1�1f3�3�3�3�34 4?4^4}4�4�4�4�5�5+6�9):Y:^:j:=#=B=a=�=$>_>�> � (   000%010c0�0�0�0,>�>�>�>�>�>   �    2�2�233(3�8w=W?   � h   �01�1�1�1�1�1�1�1�1�1222d2�2$3v3�3,4=6�9�9::$:6:V:l:�:�:�:�:�:;i;v;�;�;�;�;�;�;�;�;�;j<   �     +0�0�1�2�4�4�4�9�9???   � $   1�1225�6�7�8:�;�=�>�?   � `   �0�1�19'9E9u9�9�9:5:e:�:�:�:d;�;�<�<�<5=d=�=�=�=>#>:>C>Q>g>�>�>�>�>W?p?y?�?�?�?�?�?�? � �   0%050>0a0i0
1�1�1�2�3�3�3�34\4�4�4�4�455515C5U5g5y5�5�5�5�5�5�5�566+6=6O6a6s6�6�6�6�6�677.767�7�7�7�7 888�8�8�8
9L9P9T9X9\9`9d9h9l9p9t9�9�9�9�9�9�9�9�9�9�9�9�9�9(:,:0:4:X:\:<<'<0<n<u<X=\=`=d=h=l=p=t=x=>>f>�>�?   �   00]0{0�0�0�01�1�12,282A2�23�647p7y7�7�7�7�7�7�8�8�8�8�8�8�8�89/9<9E9�9�9�9�9:6:a:�:�:�:�:�:o;�<�<�<�<�<�<�<�<==9=L=U=�=�=�=�=�=#>+>6>A>I>�?�?�?�?    �   000"0(060>0�0�0�011"1+101E1T1c1r1�1�1 22222222303O3T3c3t3�3�3�3�3�3�3�3$4(4,4044484<4@4D4H4�4�4�4	55%5.5a5j5x5}5�5�5�5�5666p6}6�6�6�6�6�7Z8�8�8�8�8�8�8�8�8�89�9�9::!:):q;L>     "0101>1K1Z1c1|1�1�1�1�1�1�1�1�1�1x2�2�2�2�2�2�2@3`3h3n3�3�344B4M4a4l4t4�4�4�4�4�4�4�4�45$5U5�5�5�5�5>6I6`6�6�6�6�6�6�658>8c8n8�8�8�8�8�8�89!9*9M9T9a9l9�9�9�9�9�9�9:r:�:�:�:�:�:�:�: ;$;(;,;0;4;8;<;@;D;H;L;P;�;�;�;�;�;�;�;G>�>�>�>�>???H?O?�?�?�?�?�?�? 0 �   000-050T0\0c0�0�0�0�011'10151�1�1�1�1�1�1�1�1�1�1�1�1�1 2G3^3l3u3�3�3�3�3�3494�4�4�45�6�6�67	77!7E7�7�7�7t8�8�8�899%9R9�9�9�9�9�9�9�9:::J:X:a:�:�:�:;#;6;E;M;�;�;�;"<k<t<�<"=t=x=|=�=�=�=5?A?V?�?�?�?�?�? @ �   g0�0�0�0�132�3�3�3�3�3�344/4;4I4R4Y4f4o4�4�4M5d5�5�5�56$656]6t6}6�6�6�6�6�6�6�6�6777(71767H7]7l7u7�7�7�78&838u8�8�8�8�8�9�9�9�9:#:=:J:R:W:�:	<@<P<u<�<S=�=�=$>(>,>0>4>8><>@>D>H>�>�>�>�>�>   P �   0*0K0T0Z0b0k0�0�0�0�0�0�0%1�1�1�1�1�1�1I2�2�2�2�2�23n3�3�3�3�3�3�3�35�5�5�5�566}6�6�6�6�6�6�6�6�6�6�6�6�6777"7O7X7�7�7�7�7�7�7�7�7i9r9|9�9�9�9�9�9+<9<B<Q<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<=====t=x=|=�=�=�=�=�=�= ` �   50N0W0\0�011'1�1�1�122T2a2i2{2�2�2�2�2�2�3�3�3�3�3�34 4)454>4C4r4w4�4�4�4�4�4�4�4�4525?5n5{5�5�5�5�566�6v:�:�:�:�:�:�:�:�:�:	;�=�=�=@>p>�>�>�>P?�?�? p d   �1�1�1�1�1�13282A2k2p2u2�2�2�2333R3W3`3�3�3�3g5�6�8�;�;�;�;�>�>�>�>�>�> ???�?�?�?�?�?�? � X   �0�0"2d2h2l2p2t2x2|2�2
5C5H5M5P6378B9G9L9�9�9�9l:q:v:�;�;�;p<u<z<�<�<�<�>`?e?j? � <   U0�0�0'13(3u3~3 4d4i4n4:6�68	8V8%9+9::�:t;�;�=   � p   �041�3�34
424�45g6�6�6n7w7E8_8�8�8�9�9�9O:T:]:�:�:�:;8;v<{<�<�<�<�<===[=`=l=�=�=�=�=�=�=)>.>3>�>�> � x   
111B1G1L1�1�1�1�1�1�1+50595c5h5m5�5�5�5�5�5�5@;E;K;R;�;<<<o<t<}<�<�<�<:=X=�>�>�>�>�>?/?4?9?{?�?�?�?�?�?   � �   000I0N0S0�0�0=2B2G2(3-393f3k3p3�3�354:4F4v4{4�4~5�5�5�5�5�5�5y7�7�7�7�78'8U8w8�8�8939S9�:�:�:�;�<s=x=�=>>!>�?�?   � �   0A0p0�0�0
1-1O1�1�1�1�1�1�1�1(2,2024282<2@2D2H2L2�6�6�6�67$7)7b7g7p7�7�7�7:9?9H9r9w9|9�9�9�9�9�9�9
<="=.=^=c=h=�= >B>T>�>�>�>�>�>�>C?H?T?�?�?�?   � �   �014292E2u2z22!3&323b3g3l3�3{4�4�4�4�4�4�5�5�6�6�6�6�6�6888H8M8R8�9�9�9�9�9:;;%;U;Z;_;!<(<�=�=6>;>G>w>|>�>l?q?}?�?�?�?   � �   �0�0�0�0�01�1�1�1-22272$3)353e3j3o3Z4_4k4�4�4�45N6S6_6�6�6�6�7�7�7�7�7�7I8�8�9�9�9�9�9�9�:�:�:;;;�;�;�;�;�;�;�<�<�<,=1=6=>>%>U>Z>_>?�?�?�?     �   000B0G0S0�0�0)101p1w1 333A3F3K364;4G4w4|4�4`5e5q5�5�5�5�6�6�6�6�6�6�7�7�78889	99E9J9O9":':3:c:h:m:X;];i;�;�;�;�<�<�<�<�<�<�=�=�=�= >>�>�>�>?? ?  �   000L0Q0V0�5�5666;6@6�6*8/8;8k8p8u8�8�8�8�8�8�8�8�8�8�8�8 999 9$9(9,909d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9        Z?   0 �   00$0T0Y0^0�0�081J1�1�1�1�1�1�192>2J2z22�2?3u3�3�3�3 44
4X4�4�451565;566`7g7�8�8�9�:H;<<<G<L<Q<Y=>>O>V>�>�>   @ \   �5�5�5�5�56X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7e?n? P |   g0p0�0�0�0�0�0*1/181b1g1l1�3�3�3�3�3�3�4�4�4�4�4�4�5�5�5�5�5(6-626�;�;�;�<�<�<�<�<�<"='=3=`=e=j=�=�=�=�>�>�>�>�?�?�? ` �   I0N0Z0�0�0�0�0�0�0#1(1-1�1�1�1F2K2]2�2�2�2�2�2�2$3)323\3a3f364;4M4T5r5�5�5�566!6I8Q8�8�8�8
999B9G9L9�;�;�<�<�=�=#>+>�>�>�>�>Q?Y?�?�?�?�?�?�? p t   -020>0k0p0u052>2F2M2s2y2~2:6M7R7^7�7�7�7�7�7878<8A8�9�9�:�:�:*;/;4;�;�;�;<<!<o<E=L=^>c>o>�>�>�>�?�?�?�?   � �   00m1r1~1�1�1�1�2�2�2333�3�3K5R5�5�5�56!6&677$7T7Y7^7�8�8�8#9(9-9::+:[:`:e:�:<<<M<R<W<D=I=U=�=�=�=>�>~?�?�?�?�?�?   � �   �0�0�0�0�01�1�1�1�1�1�1�2�2�2333�344@4E4J4�4�5�5�5�5�5�5-626>6�6�677[7b7�8�893989=9*:/:;:k:p:u:T;Y;e;�;�;�;�<�<�<�<�<�<�=�=�=>
>>�>??=?B?G? � �   00+0[0`0e0R1W1c1�1�1�1~2�2�2�2�2�2�3�3�3�3�34�4�4�4555	666J6O6T6�;�;<3<8<=<�<>>>D>I>N>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?�?�?�?�?�?�?�? �    �?   � `   �0�0�0�0�0�0\1a1m1�1�1�1d2�2�2�2�2%3*3/3}3*414�5�5�6�689�9�:�:�:�:�:�:�;�<�<�<�<==   � h   84=4I4y4~4�4�4�4�4�4�4�4�4�4�4�4 5555$5(5,50545h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5=x=�=�=�=�>�>   � (   �0�0�011'1Q1V1[1G7�:�:�:7<�<   � X   �1�12*4�4�4�45!5&5�5�6�6#8*8	99�=�= >>>>>>>> >$>(>,>0>4>t>x>|>�>�>�>     ,   �13$3)3.3{3�3�3�3�3�3�3�344!4&4"=  h   l23-363656:6?6�6K8�:�:�:�:$;);.;g;l;x;�;�;�;�;�;�;)<.<3</=4===g=l=q=�=�=�=�=�=�=B>G>P>z>>�>     �   11)202�2�2�3�3�34@4E4N4�4�4�4�4�4�4�4#5(5-5n5s5|5�5�5�5�5"6'606i7n7z7�7�7�7�7>8C8O8|8�8�8�8�8�8�8a9f9o9�9�9�9�9�9::6:;:@:f:�:�:�:�:�:�:;?;D;M;h<�<="=A=a={=�=�=�=�=>,>M>g>�>V?e?�?�?�?�?�?�? 0 X   T0Y0b0�0�0�0�5�5E6[6�6�67@7n7�7�7�7�78
84898>8.9V9g9�9�9�9�9�9�9`:e:n:�:�:�:   @ d   001+1.3W3o3�3�4�4�4�4�45J5O5X5�5�5�5�5�5�5666�7�7�7�78	8K8P8Y8�8�8�8===�>�>�>0?<? P L   �0f2w2�2�2�2333p3u3~3�3�3�3!909J9�9�9U:k:e;{;�=�=�=�=> >%>?,?   ` �   x0}0�0�0�0�01!1*1Z1_1h1�1�1�1�1�1�122.242D2P2]2n2t2�2�2�2�2�2Q3^3y3�3�3'4[4�4�4�45�6D7m7r7w78o88�8R9W9`9�9�9�9�9�9�9:::e:j:s:�:�:�: p L   G0�0�0�0�0�0�0�1�1�2�3�34-42474�5�6W8�8�9�9�9�9�9�9z:�;�;�<�<�=�=   � �   �2�2�2�2�2�2�2�2�2�2�2�2�2 333H3L3P3�3�3�3�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�677777 7&7,72787>7D7J7P7V7\7b7h7n7t7z7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78
8888"8(8.848:8@8F8L8R8X8^8d8j8p8v8|8�8�8�8�8�8�8 �    E?u?�?�? � �   0U0�0�01:1S1z1�1�1�12=2f2�2�2
3:3j3�3�3�3U4�4�4�465f5�56�6�677�7�78+8C8[8s8�8�849t9�9�94:t:�:2;r;�;�;4<t<�<J=�=�=
>:>j>�>�>�>*?Z?�?�?�?   � �   0J0z0�0�0
1:1j1�1�1�1*2Z2�2�2�23J3z3�3�3
4:4j4�4�4�4*5Z5�5�5�56J6z6�6�6
7:7j7�7�7�7*8Z8�8�8�89J9z9�9�9*:Z:�:�:�:;B;r;�;E<v<�<�<&=S=�=�=I>v>�>�>&?S?�?�?�?   � t   0V0�0�0�061f1�1�12F2�2�2�2&3f3�3�34F4v4�4�4&5V5�5�5666v6�6�67V7�7�758�89�9�9�9?:�:)<>�>�>?O?�?�?�?   � �   0o0�0�01&1A1\1w1�1�1�1�1�1242a2�2�23!3<3W3r3�3�3�3�3�34A4�45J5z5H6H7�7�748t8�8�849t9�9�94:�:�:$;d;�;�;$<d<�<
=:=j=�=�=�=*>Z>�>�><?�?�?   �   20|0�0$1t1�1N2�2j3�3�3
4:4j4�4�4�4*5Z5�5�5�56J6�6�6�6737�7�78&8f8�8�89F9v9�9�9&:V:�:�:i<�<"=Z=s=�=�=�=�=�=>>H>�>�>�?    0   $0d0�0�0�0*1l1�12d2�223j3�3�3�3�3
4:4j4   X   o7�78_8�8�8�8�8949T9t9�9�9�9�9:4:T:t:�:�:�:�:;4;T;t;�;�;�;�;<4<T<t<�<�<�<   @ �   111111 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�2�2�2�2�2�2�2�3�3�3�3�3�3�3�3�3�3�3�3 4444444 4(4,44484@4D4L4P4X4\4`4h4l4t4x4�4�4�4�4�7�7�7�7�:�:�; P $  (0,0004080<0@0D0H0L0D1H1L1h1l1p1t1|1�1�1�1�1�1�1�1�1�1 2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�233333 3$3034383D3H3L3T3X3\3`3d3h3l3�3�3�3�3�3�3�3�3�3�3�3�3�3�34444 4�4�4�4�4�4 55555555 5$5(5,5054585H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�:�:�:�:�:�:�:�:�:�:�: ` �   $0(0�0�0�0�0�0�0�0�2�2�2�2�2�2 3$3�3�3�3�3 444$404<4H4T4`4l4x4@5L5X5d5p5|5�5�5�5�5�5�5�5�5�5`8d8h8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99   p @   0$0(0,0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01111$1,141<1D1L1T1\1d1l1t1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222$2,242<2D2L2T2\2d2l2t2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3t3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�34444$4,444<4D4L4T4\4d4l4t4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�45555$5,545<5 � �  P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�2 33333333 3$3(3,30343D3H3L3P3T3X3\3`3d3h3l3p3�3�3�3�3�3�3�3�3�3�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<$<(<,<0<4<8<<<H<L<P<T<X<\<d<h<l<p<t<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=0=@=D=H=L=P=T=X=\=`=d=h=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>$>(>,>0>4>8><>H>L>P>T>X>\>`>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????(?,?0?4?8?<?@?D?H?L?P?T?X?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�? � �   �=�=�=�=�=�=�=>>>>> >$>0>4>8><>@>D>L>P>T>X>\>`>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????(?,?0?4?8?<?@?D?H?L?P?\?`?d?h?l?   � $   �5�5�6�6�6�6�6�6 777777 �     1$1(1X9\9`9d9h9 �    �>�> ?   �    0000  �  X1`1h1p1x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 3333 3(30383@3H3P3X3`3h3p3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5(50585@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6h6p6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 8888 8(80888@8H8P8X8`8h8p8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89999$9,949<9D9L9T9\9d9l9t9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9::::$:,:4:<:D:L:T:\:d:l:t:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;$;,;4;<;D;L;T;\;d;l;t;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<<$<,<4<<<D<L<T<\<d<l<t<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====$=,=4=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\?d?l?t?|?�?�?�?       >$>(>,>0>4> 0 @   55555,747<7D7L7T7\7d7l7t7|7�7�7�7�7�7�7�7�7�7�7�7�7 `    �:�:�:�:@<D<H<   p ,   8=@=D=H=L=P=T=X=\=`=d=h=l=p=t=x=|=   �    �2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4?? ?$?,?0?4?8?@?D?H?L?T?X?\?`?h?l?p?t?|?�?�?�?   � �   h3t3�3�3�3�3�3�3�3�3�3�3�3444(444@4L4X4d4p4|4�4�4�4�4�4�4�4�4�4�4 555$505<5H5T5`5l5x5�5�5�5�5�5�5�5�5�5�5�566 6,686D6P6\6h6   � 8   00<0H0T0`0l0x0�0�0�0�0�0�0�0�0�0�0�011 1,181     �   t2(<@<X<`<t<x<�<�<�<�<�<�<�<�<�<==(=0=4=<=T=`=x=�=�=�=�=�=�=�=�=�=�= >>0>4>H>P>X>p>�>�>�>�>�>�>�>�>�>�>�>??(?@?X?\?p?x?|?�?�?�?�?�?�?�?�?�?�?�?  �  0 0$080@0D0L0d0|0�0�0�0�0�0�0�0�0 11110141H1P1T1X1`1x1�1�1�1�1�1�1�1�1�1�122222$2<2T2X2l2t2|2�2�2�2�2�2�2�2�2�233$3,3034383@3X3p3t3�3�3�3�3�3�3�3�3�3�3�3�34,404D4L4P4T4\4t4�4�4�4�4�4�4�4�4�4�4�4�4555 5$5,5D5\5`5t5|5�5�5�5�5�5�5�5�5�5�5�56,606D6L6T6l6�6�6�6�6�6�6�6�6�6�6 77 787<7P7X7`7x7�7�7�7�7�7�7�7�7 8888,8D8H8\8d8h8p8�8�8�8�8�8�8�8�8�8 999 9$9,9D9\9`9t9|9�9�9�9�9�9�9�9�9�9�9�9:: :4:<:@:D:L:d:|:�:�:�:�:�:�:�:�:�:�:�: ;; ;8;<;P;X;\;`;h;�;�;�;�;�;�;�;�;�;�;�;<<< <(<@<X<\<p<x<|<�<�<�<�<�<�<�<�<�<�<�<== =4=<=@=D=H=P=h=�=�=�=�=�=�=�=�=�=�=�=�=>>>>>0>H>L>`>h>l>p>x>�>�>�>�>�>�>�>�>�>?? ?(?,?0?8?P?h?l?�?�?�?�?�?�?�?�?�?�?�?�?�?     �  0(0,0@0H0L0P0X0p0�0�0�0�0�0�0�0�0�0�0 1111101H1L1`1h1l1p1t1|1�1�1�1�1�1�1�1�1�122$2,20242<2T2l2p2�2�2�2�2�2�2�2�2�2�2�23333$3(3<3D3H3L3P3T3`3x3�3�3�3�3�3�3�3�3�3�3�34444$4<4T4X4l4p4�4�4�4�4�4�4�4�4�4�4�4�4�45,505D5L5P5T5\5t5�5�5�5�5�5�5�5�5�5�5�56666 686P6T6h6p6t6x6�6�6�6�6�6�6�6�6�6�6�677(7@7H7L7P7T7h7l7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88 888<8P8X8\8`8h8�8�8�8�8�8�8�8�8�8�8�899(9094989<9D9\9t9x9�9�9�9�9�9�9�9�9�9�9�9�9::4:8:L:T:X:\:`:d:p:�:�:�:�:�:�:�:�:�:�:;;;;;;(;@;X;\;p;x;|;�;�;�;�;�;�;�;�;�;�;�;<< <4<8<L<P<d<l<p<x<�<�<�<�<�<�<�<�<===$=(=,=4=L=d=h=|=�=�=�=�=�=�=�=�=�= >>>0>8>@>X>p>t>�>�>�>�>�>�>�>�>�>�>�>?(?,?@?H?L?T?l?�?�?�?�?�?�?�?�?�?�? 0 \   000$0333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6$949`9h9�9�9�9�9�9�9 :D:P:X:�:�:�:�:�:;;;@;d;p;x;�;�;�;�; <$<0<8<X<`<l<p<|<�<�<�<�<�<�<�<�<�<�<�< == =,=@=L=T=`=d=p=�=�=�=�=�=�=�=�=�=�=�=�=�=>>0><>D>P>T>X>d>x>�>�>�>�>�>�>�>�>�>�>�>�>�>???(?,?8?L?X?`?l?p?t?�?�?�?�?�?�? @ �   0000<0`0l0�0�0�0�0�0�01181@1L1x1�1�1�1�1�1�1�1�1222 2H2T2|2�2�2�2�2�2�2�2�23,383\3h3�3�3�3�3�3�34$404X4`4h4p4|4�4�4�4�4�4�4�4 5(505<5d5p5�5�5�5�5�5�5�5�56$6,646@6h6t6�6�6�6�6�6�6787D7L7l7x7�7�7�7�7�7 8888 8(80888@8H8P8l8�8�8�8�8�8�8�8�8�8�8�8�8�89949@9d9l9t9�9�9�9�9�9�9�9:(:L:T:\:h:�:�:�:�:�:�:;;4;@;d;p;�;�;�;�;�; <$<0<T<`<�<�<�<�<�<�<�<�<�<�<�<==H=P=t=�=�=�=�=�=�=�=> >(>4>\>h>�>�>�>�>�>�>�>??@?`?h?p?x?�?�?�?�?�?�?�? P �   0,0P0\0�0�0�0�0�0�0�01$1,141@1h1p1x1�1�1�1�1�1�1�1 2(242X2`2l2�2�2�2�2�2�2�2�2�23,383\3h3�3�3�3�3�3�34404<4`4l4�4�4�4�4�4�4�4�4�4 5(545X5d5�5�5�5�5�5�5�56,646<6H6p6|6�6�6�6�6�67777$7,747<7D7L7T7\7d7l7t7|7�7�7�7�7�7�7888$8L8T8`8�8�8�8�8�8�8�8 9999 9(90989@9H9P9X9p9|9�9�9�9�9:,:8:@:`:h:p:|:�:�:�:�:�:�:;$;H;T;x;�;�;�;�;�;�;�;<(<L<X<|<�<�<�<�<�<==<=H=l=x=�=�=�=�=�=�=>4><>D>L>T>d>p>�>�>�>�>�> ?$?0?T?`?�?�?�?�?�?�?�? ` �   000<0D0L0T0`0�0�0�0�0�0�0�01,141@1h1p1x1�1�1�1�1�1�1�1 2202<2`2h2p2|2�2�2�2�23343@3h3�3�3�3�3�3�3�3�3�3�34,484\4d4l4x4�4�4�4�4 5555D5P5t5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6|6�6�6�6�6�6�6�6 7(747\7d7p7�7�7�7�7�7�7�7�7�7�78888$8,8D8P8t8�8�8�8�8�89949@9h9�9�9�9�9�9�9�9�9�9�9�9�9(:0:T:h:�:�:�:�:�:�:�:;(;T;x;�;�;�;�;�;�;�;�; <(<0<<<d<p<�<�<�<�<�<�<=4=@=H=h=t=�=�=�=�=�=>(>4>X>d>�>�>�>�>�>�>�>??8?@?L?t?�?�?�?�?�? p �  0040@0d0p0�0�0�0�0�0 1$101T1`1�1�1�1�1�1�1282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2�23343@3d3p3�3�3�3�3�3�3�3�3�3�3 444(4T4t4|4�4�4�4�4�4�4�4�4�455$5,545D5L5T5`5�5�5�5�5�5�5�56,686\6h6�6�6�6�6�6�6 7747T7\7d7l7t7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�78888D8h8p8x8�8�8�8�8�8�8�8(9H9P9X9`9h9p9x9�9�9�9�9�9�9�9�9�9�9 ::0:<:h:�:�:�:�:�:�:�:;;4;<;D;P;x;�;�;�;�;�;�;�;$<H<T<\<|<�<�<�<�<�<==<=H=l=x=�=�=�=�=�=�=�=>(>L>T>`>�>�>�>�>�>�>?$?L?l?t?|?�?�?�?�?�?�?�?�? � (  080D0h0�0�0�0�01(1H1h1�1�1�1�12(2H2h2�2�2�2�2�23(3D3H3h3�3�3�3�3�3�3�3�3444@4L4T4�4�4�4�4�4�4�4�4�4505P5\5h5�5�5�5�5�5�5 6 6@6`6�6�6�6�6 7 7@7`7l7�7�7�7�7 888P8p8|8�8�8�8�8�8�8909P9p9�9�9�9�9�9::(:P:p:�:�:�:�:;0;L;P;p;|;�;�;�; < <@<L<X<�<�<�<�<=0=P=p=�=�=�=�=�= >,>8>\>h>   � x   `2h2`577 7(7,7074787<7@7D7H7L7X7\7`7d7h7l7p7t7h9�9�9�9�9�9�9�9�9�9�9�9�9::::$:,:4:<:D:L:T:\:d:l:t:|:�:|?   �   x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,202<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�243\3l3|3�3�3�3�3�3�3�344044484<4@4D4H4L4P4T4`4p4t4(5,5 <H<l<�<�<�<=(=D=d=�=�=>X>�>�>?4?\?�?�?�? � �    040h0�0�0�0�0181X1|1�1�1�12@2h2�2�2�23p3�3�3$4L4p4�4 5d5�5�5�5 6h6�6�6 7�7�7�78x8�8D9l9�9�9 :�:�:�: ;h;�;�;<�<�<=4=`=�=,>P>|>�>�>�>�>?4?X?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              